�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X
   firstBloodq0X
   firstTowerq1X   firstInhibitorq2X
   firstBaronq3X   firstDragonq4X   firstRiftHeraldq5etq6bX   n_features_in_q7KX
   n_outputs_q8KX   classes_q9h"h#K �q:h%�q;Rq<(KK�q=h)X   i8q>���q?Rq@(KX   <qANNNJ����J����K tqBb�C              qCtqDbX
   n_classes_qEKX   base_estimator_qFhX   estimators_qG]qH(h)�qI}qJ(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h7Kh8Kh9h"h#K �qKh%�qLRqM(KK�qNh)X   f8qO���qPRqQ(KhANNNJ����J����K tqRb�C              �?qStqTbhEcnumpy.core.multiarray
scalar
qUh@C       qV�qWRqXX   max_features_qYKX   tree_qZcsklearn.tree._tree
Tree
q[Kh"h#K �q\h%�q]Rq^(KK�q_h@�C       q`tqabK�qbRqc}qd(hKX
   node_countqeM�X   nodesqfh"h#K �qgh%�qhRqi(KM��qjh)X   V56qk���qlRqm(Kh-N(X
   left_childqnX   right_childqoX   featureqpX	   thresholdqqX   impurityqrX   n_node_samplesqsX   weighted_n_node_samplesqttqu}qv(hnh)X   i8qw���qxRqy(KhANNNJ����J����K tqzbK �q{hohyK�q|hphyK�q}hqhQK�q~hrhQK �qhshyK(�q�hthQK0�q�uK8KKtq�b�Bg         :                   �?�2O����?�e           �@       �                    �?���G�t�?:          ���@       b                    �?`��̽�?�&           ��@       !                    �?�6��L�?�            �@                           �?p�9�A��?           ��@                           �?lٮq���?�           �@                            �?է����?�           ��@       	                     �?�@}`��?           �@������������������������       �zq�����?           0{@
                           �?ܧ��1�?            {@                           �?�BbΊ�?�            `y@������������������������       �8�'d���?�            0r@                           �?�nkK�?J            �\@������������������������       �ؗp�'ʸ??            �X@������������������������       �                     1@                           �?R�}e�.�?             :@������������������������       ���<b���?             7@������������������������       ��q�q�?             @                           �?�������?�            �u@                           �?z�RC'��?�            `p@������������������������       ��;V��?�             m@                           �?8^s]e�?             =@������������������������       ���H�}�?             9@������������������������       �                     @                           �?(�s���?8             U@������������������������       �xdQ�m��?6            @T@������������������������       �                     @������������������������       �                     @                           �?������?            �D@������������������������       �                     @                             �?@-�_ .�?            �B@������������������������       �                      @������������������������       � 	��p�?             =@"       Q                    �?`1KF5�?�           ��@#       >                    �?���)}o�?H           �@$       1                     �?���>h��?�           ؑ@%       ,                    �?\=�<�?�           h�@&       +                    �?�T �?|           x�@'       (                    �? 6,/��?r           ��@������������������������       �                      @)       *                    �?�$�'홸?p           �@������������������������       ��(.�9�?g           p�@������������������������       �        	             .@������������������������       �        
             0@-       0                    �?X�<ݚ�?U            �_@.       /                    �?�\��N��?L            �\@������������������������       ����Q��?C             Y@������������������������       �        	             ,@������������������������       �r�q��?	             (@2       ;                    �?i�rch�?           �z@3       8                    �?�+�Y]�?�            0y@4       7                    �?�K��G^�?�            @p@5       6                    �?p3����?�            �m@������������������������       �                     �?������������������������       �(2��R�?�            �m@������������������������       ��nkK�?             7@9       :                    �?z91$UO�?W            �a@������������������������       ��)z� ��?T            `a@������������������������       �                     @<       =                    �?�GN�z�?             6@������������������������       �z�G�z�?             $@������������������������       �      �?
             (@?       J                    �?�\�7��?j           h�@@       G                    �?���K ]�?/            ~@A       D                     �?���#�İ?*           �}@B       C                    �?�h����?�             u@������������������������       �@��8��?�             r@������������������������       �                     H@E       F                    �?����p�?T             a@������������������������       ����}<S�?H            �\@������������������������       �                     5@H       I                     �?���Q��?             $@������������������������       ����Q��?             @������������������������       �z�G�z�?             @K       P                    �?ʫe�s,�?;            �Z@L       O                    �?�D��?6            �X@M       N                     �?�^�����?2            �U@������������������������       ���2(&�?             F@������������������������       ��G��l��?             E@������������������������       �                     (@������������������������       �                     "@R       [                     �?���Q��?�             l@S       Z                    �?TV����?H            �]@T       W                    �?͍�@��?A            @[@U       V                    �?d�
��?5             V@������������������������       �z�G�z�?            �F@������������������������       �>��C��?            �E@X       Y                    �?���N8�?             5@������������������������       �                     @������������������������       ���S�ۿ?             .@������������������������       �                     "@\       a                    �?,y�xEE�?M            �Z@]       `                    �?zOW7���?E            @X@^       _                    �?��wy���?A             W@������������������������       ����Q��?            �A@������������������������       �x�}b~|�?)            �L@������������������������       �                     @������������������������       �                     $@c       �                    �?P �9�Ӿ?�           ��@d                           �?0����?�           ,�@e       v                    �?@���M�?A          ��@f       g                    �? ��!��?a           8�@������������������������       �        x            `g@h       o                    �?�ΉG���?�           }�@i       l                     �?�З�I�?5	           �@j       k                    �?�M�ݶ��?p           4�@������������������������       �@&2�y�?k           ��@������������������������       �                   ԓ@m       n                    �?����i�?�           h�@������������������������       ���
z���?�           x�@������������������������       �����|�p?9           �~@p       s                    �?Xc⢲K�?�	           �@q       r                     �?��c���?�           ,�@������������������������       �P䭺��?�           ��@������������������������       ��f��U˯?�           h�@t       u                     �?8
W��߰?"           |�@������������������������       ��T�4
�?e           ��@������������������������       �`��X�?�           0�@w       x                    �?����w�?�           ؇@������������������������       �                     @y       |                     �?��H>�6�?�           ��@z       {                    �?@O��F��?           |@������������������������       ������?p             g@������������������������       �p�����?�            �p@}       ~                    �?�]��?�            Ps@������������������������       �        :             U@������������������������       �Х-��ٹ?�             l@�       �                     �?�|Ȱw��?�           ��@�       �                    �?�V�K���?�           ȃ@�       �                    �?;�)���?l           h�@������������������������       ���ɜ|��?�            t@������������������������       ��Zc!J��?�            �m@������������������������       ��I�w�"�?,             S@�       �                    �?&�l�J�?           �z@������������������������       �:���u��?�            �l@�       �                    �?��q?���?�            �h@������������������������       �����.�?^             a@������������������������       �����5�?%            �N@�       �                    �?RSIY��?�           h�@������������������������       �        	             .@�       �                     �? ������?�           J�@�       �                    �?�q��uQ�?q           �@�       �                    �?�zq8�Y�?�           �@�       �                    �?x! ���?�           Ȅ@�       �                    �?H��].�?h           ��@������������������������       ��w��3(�?x            �g@������������������������       �Ȕ�f�?�            �w@������������������������       �ʂy��?I            @X@�       �                    �?h��@D��?           �z@�       �                    �?H鮜޹?�            @v@������������������������       �        G            @\@������������������������       �ؓ!'�s�?�            `n@������������������������       �L�w�=�?/            �Q@�       �                    �?�6�~笽?�            0p@�       �                    �? ���4�?�            �h@������������������������       �        !             H@������������������������       �(;L]n�?c            �b@������������������������       �L=�m��?&            �N@�       �                    �?�X�V	�?f           |�@�       �                    �?�r&]��?�           t�@�       �                    �? 5x ��?�            t@������������������������       �Pհ�*�?w            `g@�       �                    �?�����?W            �`@������������������������       ���`qM|�?2            �T@������������������������       �`'�J�?%            �I@�       �                    �?�J@Ww�?�           ��@������������������������       �t�F>s}�?            �y@�       �                    �?�G���?�            x@������������������������       �࿾��@�?w            `h@������������������������       ��˹�m��?{            �g@�       �                    �?Tr��V��?�             p@������������������������       �d�K��?P            @^@�       �                    �?�z�>#h�?V             a@������������������������       ��Z4���?'            �P@������������������������       �^������?/            �Q@�       �                    �?�ѩ!O�?[           C�@�       �                    �?�3�ŎL�?V
           &�@�       �                    �?T]����?g           \�@�       �                    �?�l�����?           �z@������������������������       �                      @�       �                    �?L�[$ś�?           `z@�       �                    �?H���e$�?�            �x@�       �                    �?4B���
�?�            �s@�       �                     �?6Vߡ��?~            �i@������������������������       �x��}�?F            �[@������������������������       ����̅��?8            �W@�       �                     �?��U/��?I            �\@������������������������       ����y4F�?/             S@������������������������       ��\��N��?             C@�       �                     �?^Gث3��?0            �S@������������������������       ��E��ӭ�?             B@������������������������       ���i#[�?             E@�       �                     �?`2U0*��?             9@�       �                    �?��S�ۿ?             .@������������������������       �                     @�       �                    �?ףp=
�?             $@������������������������       ������H�?             "@������������������������       �                     �?������������������������       �                     $@�       �                    �?��|����?[           �@�       �                    �? ����?�           D�@�       �                     �? �-�_��?�           �@������������������������       ��t����?�            �u@������������������������       ���c�|n�?�            �p@�       �                    �?�6�=ل�?K           �~@�       �                     �?@_�M�q�?           �w@������������������������       ���!���?�            p@������������������������       �        U            �^@�       �                     �?P�Lt�<�?I            �\@������������������������       �@	tbA@�?.            @Q@������������������������       �`Ӹ����?            �F@�       �                     �?�ѫ\Z�?�           Ԝ@�       �                    �?�/��:\�?�           �@�       �                    �?D�u���?D           ��@������������������������       ��8��8��?)            ~@������������������������       ��o�s(��?           �{@������������������������       ���	= ��?t            �e@�       �                    �?ܫ%���?�           ��@�       �                    �?�ܸb���?�            �@������������������������       �3���?�            �v@������������������������       �	��B�?�            Pq@������������������������       � 7���B�?C             [@�       �                    �?�2;�f�?�           ��@�       �                    �?��T�.��?�            `v@�       �                     �?      �?             @@������������������������       �������?
             1@������������������������       �                     .@�       �                     �? fQ gN�?�            `t@������������������������       ���:��?w            @f@������������������������       ����hg��?d            �b@�       �                     �?�Y񇒻�?            y@�       �                    �?nM`����?�            �l@�       �                    �?�<ݚ�?             "@������������������������       ����Q��?             @������������������������       �                     @�       �                    �?ҳ�wY;�?�            �k@������������������������       �=��T�?[            �a@������������������������       �l��
I��?/            @T@�       �                    �?�+��<��?s            �e@�       �                    �?\Ќ=��?>            �V@������������������������       �                     @������������������������       �ҳ�wY;�?:            @U@�       �                    �?�Je\���?5            @T@������������������������       �                     (@������������������������       ���x�5��?-            @Q@�                          �?���dNx�?	           :�@�                           �?�h)����?�           ؘ@�       �                    �?�a�2��?c            �@�       �                    �?f�ğ���?           �y@�       �                    �?�s��2��?�            �k@������������������������       ������?|            �g@������������������������       ��חF�P�?             ?@�       �                    �? E59|�?t             h@������������������������       �hA� �?T            �a@������������������������       ��O4R���?             �J@                          �?��0�=8�?a            `d@������������������������       ���a�n`�?H             _@������������������������       � ���J��?            �C@                         �?��[����?�           ��@                         �?|���V�?y           P�@������������������������       ��ܷ��?'           P}@������������������������       �|�űN�?R            @]@      
                   �?D�C]���?           �z@      	                   �?P�t��?,            @R@������������������������       �"pc�
�?            �@@������������������������       �P���Q�?             D@                         �?����н�?�            0v@������������������������       ��y��λ?�            pr@������������������������       �        '             N@      #                   �?�xbF��?           ��@                         �?^ۈ��.�?v            �f@                          �?���q��?L            �]@                         �?���H.�?              I@                         �?���y4F�?             3@������������������������       �d}h���?             ,@������������������������       �z�G�z�?             @                         �?�n`���?             ?@������������������������       ��+e�X�?             9@������������������������       �                     @                         �?bKv���?,            @Q@                         �?      �?             8@������������������������       ��	j*D�?             *@������������������������       �"pc�
�?             &@                         �?:	��ʵ�?            �F@������������������������       ��S����?             C@������������������������       �����X�?             @                          �?�b��-8�?*            �O@������������������������       �@�0�!��?             1@!      "                    �?���.�6�?"             G@������������������������       ��IєX�?             1@������������������������       � 	��p�?             =@$      +                   �?�g����?�           Ĝ@%      (                    �?To�ɔ�?)           0�@&      '                   �?�ј!["�?�            `v@������������������������       ���Н�z�?�            p@������������������������       ��5�uԞ�?J            @Y@)      *                   �?    ��?:            �@������������������������       ��'f��?�            v@������������������������       �l`N���?f            �c@,      3                   �?��ű?�?|           X�@-      0                   �?8OӨ�?�            Pu@.      /                    �?���9|�?�            �o@������������������������       �p���h�?O            @[@������������������������       ��5?,R�?`             b@1      2                    �?�eP*L��?8             V@������������������������       ��&!��?            �E@������������������������       �f.i��n�?            �F@4      7                   �?d�;lr�?�           ��@5      6                    �?k絊��?            {@������������������������       ��_�����?u             g@������������������������       ��7���?�             o@8      9                    �?҄��?|            �h@������������������������       ��c�����?=            �Z@������������������������       ���*(��??             W@;      r                   �?p>e�A�?�+          @B�@<      _                   �?��+���?�           ��@=      N                   �?��c)�Ǐ?�           ��@>      I                   �? �.�?Ƞ?�           ��@?      D                    �?`y����?W           H�@@      C                   �?��4+̰�?�            0r@A      B                   �?Ћ����?[            �d@������������������������       �                     �?������������������������       ���w#'�?Z            `d@������������������������       ��U���?S            �_@E      H                   �?��"pK�?�            `p@F      G                   �?���J��?B            �Y@������������������������       �                     &@������������������������       �p�C��?;            �V@������������������������       �        g             d@J      K                   �?�E��La�?i            �d@������������������������       �        -            �Q@L      M                    �?�a�O�?<            @X@������������������������       �@3����?              K@������������������������       �                    �E@O      X                   �?�A�Wb�?(           Z�@P      S                    �?@�Ҵ�3�?T           ��@Q      R                   �? �+��
�?�           ؇@������������������������       �        �            �k@������������������������       ��1Ai��?_           �@T      W                   �? �K �؁?r           l�@U      V                   �?����r�?�            �t@������������������������       �        %            �O@������������������������       � }�Я��?�            �p@������������������������       ���|�?�w?�           D�@Y      \                    �?`e	ؚ�?�            pu@Z      [                   �?�|�l�?T             a@������������������������       �`Ql�R�?            �G@������������������������       �        9            @V@]      ^                   �?@	tbA@�?�            �i@������������������������       ��i�y�?)            �O@������������������������       �@x�5?�?W             b@`      i                    �?�O�r���?           �@a      f                   �?�!�Wd�?�           ��@b      c                   �?jه��?h            �e@������������������������       �                     @d      e                   �?�+Ĺ+�?c            �d@������������������������       �:�&���?            �C@������������������������       ��m(']�?L            �_@g      h                   �?�#��ؒ}?P           @�@������������������������       �        3            �V@������������������������       �@Vהf��?           �|@j      o                   �?`���V>�?U           ܔ@k      l                   �?p���ڈ�?�            p@������������������������       �                     9@m      n                   �?��|6嗥?�             m@������������������������       � "��u�?             I@������������������������       �@��,B�?s            �f@p      q                   �?�䞠�l�?�           ؐ@������������������������       ����N8�?.            �O@������������������������       ������?�           ��@s      �                   �?�������?�           @�@t      �                    �?6�#rLs�?�           ��@u      �                   �?�����I�?�           4�@v      {                   �?    ���?P            �@w      z                   �?z�7�Z�?�            @r@x      y                   �?     ��?�             p@������������������������       ����|���?c            @c@������������������������       ��"U����?A            �Y@������������������������       ��E��ӭ�?             B@|                         �?�WR�<��?�            �k@}      ~                   �?R���Q�?k             d@������������������������       �r�0p�?I            �Z@������������������������       �H�ՠ&��?"             K@������������������������       ���Q��?(             N@�      �                   �?�;��?�           h�@�      �                   �?j����?�             o@������������������������       �|;�p)�?H            @^@�      �                   �?     ��?Z             `@������������������������       �����X�?)            �O@������������������������       ��	j*D�?1            @P@�      �                   �?X�XG��?�            @y@�      �                   �?�~$7q�?�             o@������������������������       ������x�?t            �h@������������������������       �d,���O�?            �I@������������������������       �(�Tw��?]            �c@�      �                   �?t�\�f�?           0�@�      �                   �?�����*�?I           �@�      �                   �?s��u�?�            �g@������������������������       ��"���r�?D            �X@�      �                   �?�û��|�??             W@������������������������       �lutee�?.            �P@������������������������       ����Q��?             9@�      �                   �?̳hD<�?�            �s@������������������������       �@K����?i            �d@�      �                   �?�@�q�a�?]            �b@������������������������       ��~8�e�?"            �I@������������������������       ����o_�?;             Y@�      �                   �?�P�� ��?�           ��@�      �                   �?4և����?&            |@�      �                   �?οH�G�?�            �u@������������������������       ��^�X�?<            @X@������������������������       ��=����?�            �o@�      �                   �?X&$�E�?>            �X@������������������������       �z�G�z�?             D@������������������������       ��m����?"            �M@�      �                   �?���"�?�             q@������������������������       ��D��?            �H@������������������������       ���^cY,�?�            �k@�      �                   �?�]�;�?�          ���@�      �                   �?xVD�Q�?Z           ��@�      �                   �?t���?�           ؖ@�      �                   �?�X���?�           ؇@������������������������       �                     �?�      �                    �?�&��i&�?�           Ї@������������������������       �X/�j�?           �z@������������������������       ��۵\L��?�            �t@�      �                   �?`�g�+�?�           ؅@������������������������       �                      @�      �                   �?�]��=�?�           ȅ@�      �                    �?��UV�?           �z@������������������������       ��̨�`<�?�            �o@������������������������       ��S����?q            `e@�      �                    �?H�S[��?�            �p@������������������������       �<G�7�5�?f            `d@������������������������       ��X�<ݺ?P             [@�      �                   �?�i�$[�?�           $�@������������������������       �        
             0@�      �                    �?���[Y��?�           �@�      �                   �?�¦�{��?2           ��@������������������������       �`��	��?           �x@�      �                   �?�*E
S�?-           �|@������������������������       �<;n,��?l             f@������������������������       �0� ��k�?�            �q@�      �                   �?��Y$�׾?           �@�      �                   �?dq�b���?           ��@������������������������       �@-�_ .�?           �{@������������������������       ���2(&�?h            @c@������������������������       �X`؄c�?            �x@�      �                   �?�� �{�?P           (�@�      �                   �?�ӛ��?�	           ��@�      �                   �?G��W�?B           V�@�      �                    �? ��]�?5           ��@������������������������       �І�^���?%           �|@������������������������       ����D�?           �|@�      �                    �?`OV$�2�?           .�@������������������������       ��:][^�?           (�@������������������������       ��x���?	           H�@�      �                   �?,[�_{�?�           ��@�      �                    �?tX�}}��?           P|@������������������������       ��ǟa���?�             k@������������������������       ��z���?�            �m@�      �                    �?�1�`jg�?}           �@������������������������       ����\=y�?�             k@������������������������       � ��Q�?�            @x@�      �                    �? �_aZ�?s           ��@�      �                   �? ���s�?�           �@������������������������       ��[|x��?�            �o@������������������������       ��g�y��?�           8�@�      �                   �?�����?�           `�@������������������������       � �#�Ѵ�?�            �r@������������������������       ���F���?8           ��@q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KM�KK�q�hQ�Bp      @s�@    ���@    ���@     �@    �'�@     4�@     ֠@     ��@     ��@     ��@     Ѓ@     H�@     ��@     H�@     h�@     `u@      k@     @k@     @s@      _@     �r@     @Z@     �g@      Y@     �[@      @     @W@      @      1@              @      3@      @      2@       @      �?     �Y@     `n@     �X@     �d@     �S@     `c@      4@      "@      0@      "@      @              @     �S@      @      S@              @      @               @     �C@              @       @     �A@               @       @      ;@     ��@     P{@     T�@     �r@     ��@     �n@     Ђ@     �\@     �@     �F@     �@      =@       @              �@      =@     ��@      =@      .@                      0@      L@     �Q@      K@      N@      D@      N@      ,@               @      $@     Pr@     �`@      r@     �\@     `l@     �@@     �i@      @@      �?             �i@      @@      6@      �?     �N@     �T@     �L@     �T@      @              @      1@       @       @      @      "@     ��@     �K@     �|@      4@     �|@      0@     �t@      @     �q@      @      H@             �_@      $@     @Z@      $@      5@              @      @       @      @      @      �?      R@     �A@      R@      :@      N@      :@      C@      @      6@      4@      (@                      "@     �V@     �`@     �P@      J@     �P@     �E@      G@      E@      B@      "@      $@     �@@      4@      �?      @              ,@      �?              "@      8@     �T@      8@     @R@      3@     @R@      ,@      5@      @      J@      @                      $@     ��@     @�@    ��@     ؀@    ���@     �i@     ��@      f@     `g@             ͽ@      f@     ��@      4@     �@      &@     h�@      &@     ԓ@             D�@      "@     8�@       @     �~@      �?     ڭ@     �c@     ܛ@      U@     �@     �N@     ��@      7@     ؟@      R@     H�@      C@      �@      A@     ��@      <@      @             І@      <@     {@      0@     �f@       @     `o@      ,@     �r@      (@      U@             �j@      (@     ��@     �t@     �y@     `k@     @v@      i@     �j@      [@     �a@     @W@      M@      2@     �s@      ]@     �e@     �L@     @a@     �M@     @X@     �C@     �D@      4@     N�@     �p@      .@             0�@     �p@     \�@     �[@      �@     �W@      �@     �J@     �@      ;@      g@      @     @v@      5@     �Q@      :@      x@      E@     u@      3@     @\@              l@      3@     �G@      7@     `n@      0@      h@      @      H@              b@      @      I@      &@     �@     �c@     H�@     �R@     �s@      "@      g@      @      `@      @     �S@      @     �H@       @     І@     �P@     0w@      D@     pv@      :@      g@      &@     �e@      .@     �e@     �T@     �U@      A@      V@     �H@      E@      9@      G@      8@     ��@     ��@     �@     Є@     ��@      u@     �o@      e@               @     �o@     �d@     �l@     �d@      j@     �[@      `@     @S@      U@      :@      F@     �I@      T@      A@      N@      0@      4@      2@      7@     �K@      $@      :@      *@      =@      8@      �?      ,@      �?      @              "@      �?       @      �?      �?              $@             ��@      e@      �@      1@     ��@      (@     `u@      @     p@      @     �~@      @     �w@       @     �o@       @     �^@             �[@      @      Q@      �?     �E@       @     t�@      c@     ��@     @U@     ��@      Q@     �{@      D@     �y@      <@     �c@      1@     h�@     �P@     (�@     �O@     �t@     �A@      o@      <@      Z@      @      {@     �t@     �g@     �d@      @      <@      @      *@              .@     `g@     `a@     �X@      T@     @V@     �M@      n@      d@      b@     @U@       @      @       @      @              @     �a@     �S@     �U@      K@     �L@      8@      X@      S@     �K@      B@              @     �K@      >@     �D@      D@              (@     �D@      <@     ܟ@     ��@      �@     ؐ@     0p@     �s@      j@     �i@      7@     �h@      2@     `e@      @      :@     @g@      @     �`@      @      J@      �?      I@     @\@      (@      \@      C@      �?     �o@     ȇ@     �`@     `|@      7@     �{@     @[@       @     @^@     0s@      F@      =@      @      ;@      C@       @     @S@     `q@      1@     `q@      N@             ܗ@      @      P@     �]@     �G@      R@      5@      =@      .@      @      &@      @      @      �?      @      9@      @      3@              @      :@     �E@      2@      @      "@      @      "@       @       @     �B@      @      @@       @      @      1@      G@      ,@      @      @     �E@      �?      0@       @      ;@     ܖ@     �w@     ��@     �h@      r@     �Q@      m@      9@      L@     �F@     �w@      `@      r@     �O@     @W@     �P@     ��@     `f@      q@     @Q@      m@      5@     @Y@       @     ``@      *@      D@      H@      :@      1@      ,@      ?@     @�@     �[@     px@     �D@     �d@      3@     @l@      6@      `@     @Q@      T@      :@     �H@     �E@     �@     ��@     �I@     V�@      9@     Ȩ@      (@      �@      &@     ��@      "@     �q@      @     �c@              �?      @     �c@      @      _@       @     @p@       @      Y@              &@       @     @V@              d@      �?     �d@             �Q@      �?      X@      �?     �J@             �E@      *@     @�@      "@     ��@      @     ��@             �k@      @     Ѐ@      @     T�@      @     pt@             �O@      @     �p@      @     8�@      @     0u@      �?     �`@      �?      G@             @V@      @     �i@       @     �N@      �?     �a@      :@     ȟ@      ,@     8�@      (@      d@              @      (@     @c@      @      @@      @     �^@       @     0�@             �V@       @     �|@      (@     ��@      @     �o@              9@      @     `l@      @     �G@       @     �f@      @     ��@      @      N@      @     ��@      �@     \�@     ��@     �@     pv@     0�@      d@     �u@      Z@     �g@     �W@     @d@      L@     �X@      C@      P@      $@      :@     �L@     `d@      B@      _@      =@     @S@      @     �G@      5@     �C@     �h@     p|@      U@     �d@      G@     �R@      C@     �V@      2@     �F@      4@     �F@     �\@      r@     �K@      h@      E@     `c@      *@      C@     �M@     @X@     p{@     ��@     �j@     pr@     �S@      \@     �E@      L@      B@      L@      :@     �D@      $@      .@     �`@     �f@     @Q@     @X@     @P@     �U@      6@      =@     �E@     �L@     @l@     �~@      c@     pr@     �\@     @m@      >@     �P@     @U@     �d@      C@     �N@       @      @@      >@      =@     @R@     �h@      *@      B@      N@     `d@     P�@    �>�@     t@     |�@      f@     �@      V@     �@              �?      V@     �@     �G@     �w@     �D@     Pr@      V@     �@               @      V@     �@      K@     @w@      ;@     �l@      ;@      b@      A@     �m@      <@     �`@      @     �Y@      b@     ��@              0@      b@     ��@     @T@     0�@     �E@     �u@      C@     �z@      *@     `d@      9@     Pp@      P@     �@     �F@     H�@      8@     @z@      5@     �`@      3@     �w@     �v@     ��@     @m@     ƭ@     �c@     �@     �J@     ��@      9@     �z@      <@      {@     �Y@     ��@     �J@     ��@      I@     ��@     �S@     ��@     �F@     �y@      1@     �h@      <@      j@     �@@     ��@      2@     �h@      .@     Pw@     �_@     ��@     �F@     ��@      4@      m@      9@     p�@     �T@     �@      ,@     �q@      Q@     ��@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q��q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheM�hfh"h#K �q�h%�q�Rq�(KM��q�hm�BXh         :                   �?$��W��?f           �@       �                    �?��U�y�?:          @��@       r                    �?^*N��?�           ĳ@       C                    �?H���E�?|
           ��@                           �?8&��[�?9           �@                           �?������?�           ��@                           �?�\]�{�?�           x�@                            �?l+�����?S           �@	       
                     �?d���W��?�           @�@������������������������       ���s����?           �{@������������������������       �����`�?�            �p@������������������������       ���|��?�            `o@                            �?��F��?c            `c@                           �? _�@�Y�?J             ]@                           �?0�)AU��?I            �\@������������������������       �@��8��?>             X@������������������������       �                     2@������������������������       �                      @                           �?8�Z$���?            �C@                           �?�S����?             C@������������������������       �д>��C�?             =@������������������������       ������H�?             "@������������������������       �                     �?                           �?      �?C             X@                            �?��� ��?@            @W@������������������������       ������?             3@������������������������       ��L���?3            �R@������������������������       �                     @       6                    �?
�\�k��?@           @�@       '                     �?�bv}9��?           8�@       &                    �?h� ��y�?�           T�@        #                    �?��<����?�           $�@!       "                    �?p��ˮ?$           0�@������������������������       ���4+̰�?i           0�@������������������������       �      �?�             r@$       %                    �?噼:��?_            `d@������������������������       �`3�a���?E            �\@������������������������       � \� ���?            �H@������������������������       �        -             S@(       1                    �?F�FE���?g           ȁ@)       .                    �?�i��D�?�            �x@*       -                    �?�>W{�U�?�            �v@+       ,                    �?��w\ud�?�            �m@������������������������       �                     @������������������������       �H�f�i��?�            @m@������������������������       �     ��?P             `@/       0                    �?�FVQ&�?            �@@������������������������       �HP�s��?             9@������������������������       �                      @2       5                    �?�|�
��?m            @e@3       4                    �?,����?]             b@������������������������       �4��?�?D             Z@������������������������       �D^��#��?            �D@������������������������       �                     9@7       >                    �?"pc�
�?)            �P@8       ;                     �?¦	^_�?             ?@9       :                    �?�t����?             1@������������������������       �z�G�z�?
             .@������������������������       �                      @<       =                    �?����X�?
             ,@������������������������       ��q�q�?             "@������������������������       �z�G�z�?             @?       B                    �?�#-���?            �A@@       A                     �? �Cc}�?             <@������������������������       �                     $@������������������������       �r�q��?	             2@������������������������       �                     @D       [                     �?���t�?C           ��@E       P                    �?Si��?X            �@F       M                    �?nIiK���?�            �m@G       J                    �?#n��?�            �j@H       I                    �?����9�?             i@������������������������       ��1��!�?U            �`@������������������������       ��� =[�?*             Q@K       L                    �?؇���X�?
             ,@������������������������       ������H�?             "@������������������������       �z�G�z�?             @N       O                    �?�C��2(�?             6@������������������������       �                     0@������������������������       ��q�q�?             @Q       T                    �?�O*_��?�            ps@R       S                    �?pe����?�            �p@������������������������       ���i���?�            �l@������������������������       �H�V�e��?             A@U       X                    �?�LQ�1	�?             G@V       W                    �?     ��?             0@������������������������       �؇���X�?             @������������������������       ��<ݚ�?             "@Y       Z                    �?ףp=
�?             >@������������������������       �ȵHPS!�?             :@������������������������       �                     @\       e                    �?��&Zf�?�           �@]       b                    �?��(��r�?�           ؄@^       _                    �?vA����?S            ``@������������������������       �                     �?`       a                    �?D������?R            @`@������������������������       ����̅��?=            �W@������������������������       �">�֕�?            �A@c       d                    �?�HV�攽?U           ��@������������������������       �HN\�
Ե?=           �~@������������������������       ��%^�?            �E@f       k                    �?�������?C            �Y@g       j                    �?��%��?            �B@h       i                    �?�KM�]�?             3@������������������������       ��8��8��?             (@������������������������       �؇���X�?             @������������������������       �                     2@l       o                    �?r٣����?+            �P@m       n                    �?և���X�?             5@������������������������       ��eP*L��?             &@������������������������       ��z�G��?             $@p       q                    �?�:�^���?            �F@������������������������       ���p\�?            �D@������������������������       �      �?             @s       �                    �?��qu�?           ��@t       �                    �?�l�R�?�           (�@u       �                    �?�g�����?t             f@v       {                     �?��cܽ��?g            `c@w       z                    �?�&!��?:            �U@x       y                    �?Ȩ�I��?             �J@������������������������       �                     @������������������������       �H.�!���?             I@������������������������       �����e��?            �@@|                           �?(���X�?-            @Q@}       ~                    �?����e��?            �@@������������������������       �                      @������������������������       ��P�*�?             ?@������������������������       �tk~X��?             B@������������������������       �                     5@�       �                    �?,�H�Q<�?T           P@�       �                    �?�������?W            ``@�       �                     �? �q�q�?             8@������������������������       �                     @������������������������       ��X�<ݺ?             2@�       �                    �?ް� ��?G            �Z@�       �                     �?�q��/��?@            �X@������������������������       ����y4F�?             C@������������������������       ���S�ۿ?(             N@�       �                     �?�q�q�?             "@������������������������       ����Q��?             @������������������������       �                     @�       �                     �?Ȥ4"��?�             w@�       �                    �?`�q�0ܴ?>            �W@������������������������       ��g�y��?=            @W@������������������������       �                     �?�       �                    �?���.�6�?�            @q@������������������������       ������?�            �p@������������������������       �      �?              @�       �                    �? 5x ��?>            �Z@�       �                     �?�C��2(�?             6@�       �                    �?z�G�z�?             $@������������������������       ��q�q�?             @������������������������       �                     @������������������������       �        	             (@�       �                     �?`��>�ϗ?/            @U@�       �                    �?��<b�ƥ?             G@������������������������       �                     2@������������������������       �h�����?             <@������������������������       �                    �C@�       �                    �?��d��?�-          @ �@�       �                    �?�IQu`�?f           ��@�       �                    �?�s���?�          ���@�       �                    �?XE^f��?6           ��@������������������������       �        U            @`@�       �                     �?0G���ջ?�
           �@�       �                    �?`��Ȝ��?           B�@�       �                    �?WFw:�?4           ��@������������������������       �@c����?O           @�@������������������������       �pľ��l�?�           0�@������������������������       ���`��?�            Pt@�       �                    �?(��g3	�?�           ��@�       �                    �?��'cy�?K           ��@������������������������       �`��'2��?�           (�@������������������������       ��0Vq�?�           ��@������������������������       �ڲ�-���?�            �i@�       �                     �?��i�~�?�           �@�       �                    �?�c��Jj�?L           d�@�       �                    �?�U��Ԡ?~           ֧@�       �                    �?@��+S��?R           �@������������������������       �        �           (�@�       �                    �?�l��8��?W           ��@������������������������       �                     @������������������������       ���P���?S           �@�       �                    �?@:��JU�?,           @~@�       �                    �?`�LVXz�?u            �h@������������������������       �                     @������������������������       ��q�q�?q             h@������������������������       ��w�uz
�?�            �q@�       �                    �?nzMv��?�            pt@������������������������       ��R�Z��?�             p@������������������������       ���<b���?+            @Q@�       �                    �?(�0����?5           �@�       �                    �?(q�|�?�           �@������������������������       �                     ,@�       �                    �?(SH�]��?�           ��@�       �                    �?�q4t��?�           0�@������������������������       ��}3+lڎ?A           x�@������������������������       �ԓ���?�           �@�       �                    �? Um*n�?�            r@������������������������       ��q�q�?>             X@������������������������       ����|$ö?}             h@�       �                    �?     ��?�             h@������������������������       �pܹn��?b            �a@������������������������       ���[�8��?            �I@�       �                     �?��@�	�?�           ��@�       �                    �?(�0**�?P           T�@�       �                    �?��O5�?�           Ԑ@������������������������       �                      @�       �                    �?��/�V�?�           ��@�       �                    �?x�����??           ��@�       �                    �?�+�h��?�            Pq@������������������������       ���v$���?p            �f@������������������������       �        =            �W@�       �                    �? J�'.��?�           ��@������������������������       �p�u$v��?�            �v@������������������������       �Hm_!'1�?�            �n@�       �                    �?���"͏�?r             g@������������������������       �$f����?B            @]@������������������������       �H�V�e��?0             Q@�       �                    �?�h����?�             l@�       �                    �?��즟E�?x            �e@������������������������       �                     E@������������������������       �@M^l���?]            �`@������������������������       ����c�H�?#            �H@�       �                    �?�t
���?_           �@������������������������       �                      @�       �                    �?L��a��?]           �@�       �                    �?�z�oe�?�           ��@�       �                    �?��j���?�           ��@�       �                    �?��&��\�?b           ؀@������������������������       ���$����?s            �e@������������������������       �ة�!�J�?�            �v@������������������������       ��z�G��?]            �b@�       �                    �?�L���?�            �t@�       �                    �?�@�+�?�            �q@������������������������       � �)���?1            @T@������������������������       �8?W���?{             i@������������������������       ���x_F-�?#            �I@�       �                    �?�+ت�M�?�            �s@�       �                    �?x�U���?�            �m@������������������������       �lGts��?$            �K@������������������������       ����.�6�?x             g@������������������������       �����X�?3            @S@�       #                   �?<1�K���?-           1�@�                          �?L�Og���?�           �@�                          �?�6L"�?�           ��@�       �                     �?�2
�ޗ?�           ��@�       �                    �?�2�T�I�?�           ��@�       �                    �? qzu��?�           ��@������������������������       � �?����?�            pw@������������������������       �@�?B�?�            �q@������������������������       ��J�T�?,            �Q@�                           �?��E>W]�?            �|@�       �                    �?@>�Q�?            z@������������������������       �����e��?�            �p@������������������������       � i�*$Ŋ?a             c@������������������������       �`���i��?             F@      	                   �?@�?1X�?           �|@                         �?�����?�            �u@                          �?��d�?�             o@������������������������       ��t:ɨ�?Q            �`@������������������������       �XB���?J             ]@                          �?T��,��?:            @Y@������������������������       �                    �F@������������������������       ��h����?             L@
                          �?����q�?D            @[@������������������������       �                     C@������������������������       ��J�T�?)            �Q@                          �?	W�FN�?�           ��@                         �?W��Z�?I           �@                         �?��9���?�           ��@������������������������       �|T(W�j�?:           �~@������������������������       � Ϸ�~�?�             r@                         �?��{�B�?a           ��@                         �?��0_�,�?g           ȁ@������������������������       ��gߒm��?           P{@������������������������       ��5[|/��?Z            �`@                         �?������?�            �w@������������������������       ��#-���?w            �e@������������������������       ��P�I[��?�            �i@                         �?�|���?�           Ж@                         �?�NW���?�           0�@                         �?E2X�?�           �@������������������������       ���`ۻ��?�            �w@������������������������       ��{��?�            �p@������������������������       ��C��2(�?F            �X@                          �?������?�           p�@������������������������       �H�z���?�             t@!      "                   �?H"Б$�?�            �x@������������������������       �\#r��?Q            �^@������������������������       ��θV�?�            @q@$      /                    �?H4���?S           (�@%      *                   �?��U\�?�?�           ��@&      '                   �?�!�,�E�?           `{@������������������������       ����Q��?�             i@(      )                   �?F��2<��?�            �m@������������������������       �2ox��?`            �c@������������������������       �,ZYN(��?8            @T@+      ,                   �?n���6�?�            �q@������������������������       �.T�߸��?J             _@-      .                   �?�r�K��?Z            `d@������������������������       ��lg����?            �E@������������������������       ����Q��?D             ^@0      5                   �?J�w�*��?�           ��@1      2                   �?�5g����?�            pt@������������������������       �R��	P�?Z            �`@3      4                   �?�q�q�?v             h@������������������������       ��q�q�?F             ^@������������������������       ��q�q�?0             R@6      7                   �?�Ճ �?�            �r@������������������������       �.���ڨ�?g            �c@8      9                   �?�ƥ���?[            �a@������������������������       �\�����?!            �K@������������������������       � 9�����?:             V@;      �                   �?�+�����?�+          �H�@<      c                   �?��#�(�?          ��@=      T                   �?`�M#.�?W           f�@>      I                   �?@tM�?k           ��@?      D                    �?�f�¦ζ?�            t@@      C                   �?Pq�����?i            @e@A      B                   �?      �?Q             `@������������������������       �                     @������������������������       �`Jj��?O             _@������������������������       �                     E@E      H                   �?���	���?b            �b@F      G                   �?���>4ֵ?K             \@������������������������       �                      @������������������������       ���s�n�?F             Z@������������������������       ��7��?            �C@J      O                    �?�Q�A�?�           ؄@K      N                   �?@v�����?�             n@L      M                   �?���ʄ?s            �h@������������������������       �                     4@������������������������       � J���#�?h             f@������������������������       �                     F@P      Q                   �?����P��?           �z@������������������������       �        1            �Q@R      S                   �? ���,\�?�            @v@������������������������       �`�LVXz�?�            �r@������������������������       ����#�İ?'            �M@U      \                   �?@Q�g�9�?�           ��@V      Y                   �?�Qy©��?           0�@W      X                    �?�]���?�            �u@������������������������       � �)���?g            @d@������������������������       ��~��?n            �f@Z      [                    �? nT�\|?@           ��@������������������������       ��V=��|?y           8�@������������������������       � �f|�|?�           ��@]      `                   �?`ִ�[�?�            �s@^      _                    �?���J��?B            �Y@������������������������       � �q�q�?#             H@������������������������       �                     K@a      b                    �? j'����?�             k@������������������������       �        ?            �U@������������������������       � ����?V            @`@d      �                   �?      �?�           ��@e      t                   �?�
$CKr�?+           X�@f      m                   �?�s��ǝ�?�           8�@g      j                   �?R� �0�?           px@h      i                    �?ھ�l��?�            �m@������������������������       �������?^            �a@������������������������       ��fSO��?@            �X@k      l                    �?���=A�?n             c@������������������������       �VP��g��??             W@������������������������       ��0u��A�?/             N@n      q                   �?����q�?�             v@o      p                    �?�q�/;q�?�            �j@������������������������       ���VT4�?N            �\@������������������������       �r٣����?;            �X@r      s                    �?��<b���?P            @a@������������������������       �n�C���?3            �V@������������������������       ���E�B��?            �G@u      |                   �?|җ�rO�?F           x�@v      y                    �?<�:z]�?�            �w@w      x                   �?tݹ��B�?b            `c@������������������������       ��9�z���?>            @Y@������������������������       �������?$             K@z      {                   �?�ćo�?�            @l@������������������������       ��8�jC��?l            `f@������������������������       �p�v>��?             �G@}      �                   �?�kp��E�?X           ��@~                          �?�7���?           `}@������������������������       ���[�p�?n            �g@������������������������       �Z�K�D��?�            �q@�      �                    �?�x�(��??             W@������������������������       �������?            �F@������������������������       ���C���?"            �G@�      �                   �?���l]��?�           b�@�      �                    �?0�N�]��?P           ��@�      �                   �?@a���)�?p           d�@�      �                   �?l
�J�?8           h�@������������������������       ���5�n��?�            �x@������������������������       �x&xg�`�?:           �}@�      �                   �?��w��?8           �~@������������������������       �     '�?�             p@������������������������       ��#%�l��?�            �m@�      �                   �?�B!A�?�           ��@�      �                   �?��
O:�?%           �{@�      �                   �?P�I;l�?�            �q@������������������������       �                     @������������������������       ���� ��?�            pq@������������������������       �P5�޷�?k            �c@�      �                   �?@�?���?�           ��@������������������������       ��IєX�?&           �|@������������������������       �"��,;�?�            �l@�      �                   �?����>l�?L	           B�@�      �                    �?D�ۀ+�?�           ��@�      �                   �?�d<��_�?_           8�@������������������������       �                     @�      �                   �?DS���|�?]            �@������������������������       ��!N��:�?           `y@������������������������       �,�d�vK�?[            �a@�      �                   �?������?t           ��@�      �                   �?��?���?           �z@������������������������       �                     @������������������������       ��!ʉ�?
           `z@�      �                   �?��(�#H�?g            �d@������������������������       �                      @������������������������       ��r����?f            �d@�      �                    �?P��t�y�?y           R�@�      �                   �?�J�M��?�           �@������������������������       ��N^��M�?           ��@������������������������       �8�G�V޳?�             q@�      �                   �?0����ָ?�           ��@������������������������       ����D�޹?�           ��@������������������������       �xEہ@ô?�            0s@�      �                   �?&&#[��?�           ��@�      �                   �?N�UV��?           <�@�      �                   �?,�-�h��?�            �x@�      �                    �?��G���?`            �b@�      �                   �?���N8�?.            �O@������������������������       �z�G�z�?             >@������������������������       ����!pc�?            �@@�      �                   �?,�"���?2            @U@������������������������       �@��8��?             H@������������������������       �4�B��?            �B@�      �                    �?��r._�?�            �n@�      �                   �?>�ԛ���?S            �_@������������������������       �@	tbA@�?4            @Q@������������������������       ���o	��?             M@�      �                   �?�t����?L            �]@������������������������       ���v$���?)            �N@������������������������       �^l��[B�?#             M@�      �                    �?X8����?           (�@�      �                   �?P����?�             x@������������������������       �`���4�?g            �e@������������������������       ������?�            �j@�      �                   �?������?           0|@�      �                   �?��.N"Ҭ?^            @a@������������������������       �                     �?������������������������       ��ㄡ^�?]             a@������������������������       ��0ծ5��?�            �s@�      �                   �?(l��ڿ?�           )�@�      �                   �?�]ղ��?           T�@������������������������       �                     L@�      �                    �?��ɍ!��?�           t�@�      �                   �?�S����?1           �~@������������������������       � ��+&ɐ?P            @^@�      �                   �?�)�Db��?�            @w@������������������������       �H���I�?+            �S@������������������������       ���5�l@�?�            Pr@�      �                   �?�z�b��?�           ��@������������������������       ��)�"*�?r             e@�      �                   �?p�zk��?R           8�@������������������������       ��ʻ����?B            �Y@������������������������       ���	�?           z@�      �                    �?��Ujѡ�?�	           ��@�      �                   �?�L9ҁ�?Q           �@������������������������       ��u9'�ɂ?            {@�      �                   �?Ȉ�����?=           ��@������������������������       ��r����?W            �`@������������������������       ��nkK�?�           p�@�      �                   �?���7�?[           �@������������������������       � �h{��v?�           Ȑ@�      �                   �?`�l��l�?�           l�@������������������������       ��3��^�?~             h@������������������������       ��#>�	q�?D           h�@q�tq�bh�h"h#K �q�h%�q�Rq�(KM�KK�q�hQ�B�      @f�@    ���@    ���@     �@     L�@     <�@     :�@     \�@     h�@     Њ@     �@     ��@     ��@     �~@     0~@      ~@     �x@     �s@      l@     `k@     �e@      X@     �U@     �d@     `b@       @     �\@       @      \@       @     �W@       @      2@               @             �@@      @      @@      @      8@      @       @      �?      �?              (@      U@      (@     @T@      @      *@      @      Q@              @     Ȗ@     �q@     ��@      m@     ȏ@      W@     h�@      W@     X�@      ;@     ��@      2@     pq@      "@     �X@     @P@     �N@     �J@     �B@      (@      S@             �z@     �a@     0r@      [@     @p@     �Z@      j@      =@      @             �i@      =@     �I@     @S@      ?@       @      7@       @       @             @a@      @@     @\@      @@     �W@      $@      3@      6@      9@              (@      K@      "@      6@      @      (@      @      (@       @              @      $@      @      @      �?      @      @      @@      @      9@              $@      @      .@              @     �v@     �@     `l@     t@     @f@     �M@      f@     �C@     �d@     �B@     �Z@      :@     �L@      &@      (@       @       @      �?      @      �?       @      4@              0@       @      @     �H@     `p@     �@@      m@      :@     �i@      @      ;@      0@      >@      *@      @      @      �?      @       @      @      ;@      @      7@              @     �`@     ��@     @Y@     ��@      Q@     �O@              �?      Q@      O@      F@     �I@      8@      &@     �@@     p@      6@     p}@      &@      @@     �@@     �Q@      1@      4@      1@       @      &@      �?      @      �?              2@      0@      I@      (@      "@      @      @      @      @      @     �D@      @      C@      �?      @      a@     8�@     �`@     ��@     @W@     �T@      R@     �T@      J@      A@     �C@      ,@              @     �C@      &@      *@      4@      4@     �H@      *@      4@               @      *@      2@      @      =@      5@             �D@     �|@      3@      \@      �?      7@              @      �?      1@      2@     @V@      (@     �U@       @      >@      @      L@      @      @       @      @      @              6@     �u@      @     �V@      @     �V@      �?              2@      p@      (@      p@      @       @      @      Z@       @      4@       @       @       @      @              @              (@      �?      U@      �?     �F@              2@      �?      ;@             �C@    @d�@     ��@     r�@     `�@     ��@     �@     ��@     �o@     @`@             �@     �o@     �@     �b@     .�@     @Q@      �@       @     <�@     �N@     �n@     @T@     $�@     �Y@     ��@      J@     ��@      @     x�@     �F@     �c@      I@     �@     p@     .�@     `c@     p�@     �I@     ̣@     �@@     (�@             p�@     �@@      @             `�@     �@@      }@      2@     �h@       @      @             �g@       @     �p@      0@     �k@      Z@      e@     @V@      K@      .@     T�@     �Y@      �@     �I@      ,@             �@     �I@     ��@     �D@     X�@      @     ��@     �B@     pq@      $@     �W@      �?      g@      "@     �a@     �I@     @Y@      D@      D@      &@     Ģ@     �m@     Ē@      Y@     �@      V@       @             ��@      V@     H�@     �E@      q@      @     �f@      @     �W@             ��@      D@     `u@      4@      l@      4@     �a@     �F@     �U@      ?@      K@      ,@     �j@      (@     �e@      �?      E@             �`@      �?      C@      &@     Ē@     `a@       @             ��@     `a@     ،@     �X@     H�@      R@      �@      ;@      e@      @     pu@      8@     @Z@     �F@      s@      ;@     �p@      1@      T@      �?      g@      0@     �D@      $@     @q@      D@     �k@      2@     �H@      @     �e@      (@     �K@      6@     ��@      �@     ��@      u@     D�@      <@     T�@      ,@     x�@       @     P�@      @     0w@      @     pq@       @     @Q@       @     `|@      @     �y@      @     @p@      @     �b@      �?     �E@      �?     �{@      ,@     u@      (@     �m@      "@     �_@      @      \@      @     �X@      @     �F@             �J@      @     �Z@       @      C@             @Q@       @     ��@     @s@     ��@     �b@     ��@     �T@     �{@      H@      p@      A@     ��@     @Q@     Ȁ@      @@     �y@      9@     @_@      @     pu@     �B@      d@      .@     �f@      6@     \�@     �c@     p�@      L@     ��@     �G@     �u@      >@     @o@      1@     �V@      "@     H�@     @Y@     0p@     �N@     `v@      D@     �[@      (@      o@      <@     ��@     ��@      z@     0s@     �o@     @g@      ^@      T@     �`@     �Z@     �T@     �R@     �H@      @@     �d@     @^@     �P@     �L@     �X@      P@      ;@      0@      R@      H@     @w@     p@     `h@     �`@     �T@      J@      \@      T@     �Q@      I@      E@      >@      f@     @_@     @Y@      M@      S@     �P@      =@      :@     �G@     �D@     ��@    ���@     �@    ��@     �B@     �@      5@     8�@      .@      s@       @     @d@       @      ^@              @       @      ]@              E@      @      b@      @     �Z@               @      @     �X@       @     �B@      @     ��@      �?     �m@      �?     `h@              4@      �?     �e@              F@      @     `z@             �Q@      @     �u@      @     `r@       @     �L@      0@     ��@      (@     �@      @     0u@       @      d@      @     `f@      @     �@       @     (�@      @     Б@      @     �s@       @      Y@       @      G@              K@       @     �j@             �U@       @      `@     ��@     �@     h�@     $�@     @m@     �@     �b@     @n@     �X@     �a@     �J@     �U@      G@     �J@      I@     �Y@      ;@     @P@      7@     �B@     @U@     �p@     �K@     �c@      ?@      U@      8@     �R@      >@      [@      8@     �P@      @     �D@     0r@     `�@     �]@     pp@     �B@     �]@      7@     �S@      ,@      D@     @T@      b@     �P@      \@      ,@     �@@     �e@     Px@     �a@     �t@      D@     �b@     �Y@     �f@      ?@     �N@      (@     �@@      3@      <@      }@     ��@     �k@     ʡ@     �]@     ��@      R@     (�@     �G@      v@      9@     P|@      G@     �{@      ;@     �l@      3@      k@     �Y@     �@     �J@     0x@      B@     �n@              @      B@     `n@      1@     �a@     �H@     ��@      ;@      {@      6@     �i@     �n@     V�@     �X@     X�@      L@     �~@              @      L@     �~@     �F@     �v@      &@     ``@      E@     8�@      4@     `y@              @      4@      y@      6@      b@               @      6@     �a@     �b@     *�@     �Q@      �@      N@     ؇@      &@     Pp@     @S@     T�@      P@     ��@      *@     `r@     �}@     �@     �`@     $�@     �Q@     @t@      <@      ^@      .@      H@      @      8@      "@      8@      *@      R@      �?     �G@      (@      9@      E@     �i@      <@     �X@      �?      Q@      ;@      ?@      ,@     @Z@      �?      N@      *@     �F@      P@     (�@      E@     �u@      9@     �b@      1@     `h@      6@     �z@      @     �`@              �?      @     �`@      2@     pr@     �u@     Ѳ@      `@     T�@              L@      `@     t�@     �J@     �{@      �?      ^@      J@      t@      <@     �I@      8@     �p@     �R@     (�@       @     �d@     @R@     �{@     �F@     �L@      <@     Px@      k@     ��@     @V@     ��@       @      {@     �U@     ��@     �J@     �T@      A@     `�@     �_@     �@      @     ��@      _@     |�@      P@      `@      N@     x�@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q��q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheM�hfh"h#K �q�h%�q�Rq�(KM��q�hm�BXh         8                   �?D�].��?�e           �@       �                    �?Z�i���?:           �@                           �?\�U���?�(           (�@       	                    �?F�8����?Q           �@                            �?Pr=x)��?K           ��@                            �?� q��?�           ��@������������������������       �������?           0|@������������������������       �>��y���?�            `o@������������������������       ����I���?�            �k@
                            �?؇���X�?             @������������������������       �                      @                           �?z�G�z�?             @������������������������       �                      @������������������������       ��q�q�?             @       |                    �?|��.��?]&          �~�@       M                    �?�vg��?�!           ��@       0                    �?`=^n�?-          ���@       '                    �?p�K.B��?�           ��@       "                    �?P^QV=�?�           ؕ@                            �?�M��qĿ?Q           t�@                           �?x ����?_           ،@                           �?�q�q�?A             X@������������������������       �����ȫ�?6            �T@������������������������       �                     ,@                           �?h�� MQ�?           ؉@������������������������       ��8�G�ֹ?c            �@������������������������       ��/R���?�            �q@                           �?°	~��?�             x@                           �?��Pd�]�?�            `q@������������������������       �R���Q�?             D@������������������������       �����n�?�            �m@        !                    �?X'"7��?H             [@������������������������       �                     @������������������������       ����N8�?F            @Z@#       &                     �?(����7�?5            @V@$       %                    �?�c�����?!            �J@������������������������       �                      @������������������������       ���[�8��?             �I@������������������������       ��q�q�?             B@(       /                    �?io8�?H             ]@)       ,                     �?*
;&���?             G@*       +                    �? �Cc}�?             <@������������������������       �                     @������������������������       �H%u��?             9@-       .                    �?�<ݚ�?             2@������������������������       �                     �?������������������������       �������?             1@������������������������       �        +            �Q@1       <                     �?��NK�?_          ���@2       3                    �?@�v��ġ?(           V�@������������������������       �        \            �`@4       7                    �?����.�?�           ҵ@5       6                    �? �ձ��t?�           b�@������������������������       �@�6�Ds�?t           ̕@������������������������       �        n           ��@8       ;                    �?�V-y�U�?�           B�@9       :                    �?�j	�ڬ?5           �@������������������������       ��,���)�?�           ��@������������������������       �Pe ����?Z           T�@������������������������       ���Ú���?�            �r@=       F                    �?(�E���?7           �@>       A                    �?�ʏ��X�?!           �@?       @                    �? >��
�?�           �@������������������������       �                     7@������������������������       � q7V��?�           `�@B       C                    �? ôZC7k?�           Ȃ@������������������������       �        	             4@D       E                    �? �¯&l?z           (�@������������������������       ����1��p?:            ~@������������������������       �        @            �X@G       H                    �?��(�S�?           <�@������������������������       �                     "@I       L                    �?����n2�?           �@J       K                    �?���(�޹?�            �@������������������������       ��Va����?�           ȇ@������������������������       �0�hg���?�           x�@������������������������       ��˹�m��?}            �g@N       e                    �?�I��-�?m           
�@O       Z                    �?�Fa/���?�           ��@P       W                    �?���L��?            �x@Q       T                    �?R���2��?�            �t@R       S                     �?X閘��?�            `l@������������������������       �\�CX�?^            �a@������������������������       �Ї?��f�?6            @U@U       V                     �?r�0p�?@            �Z@������������������������       ����@��?+            �R@������������������������       �     ��?             @@X       Y                     �?V��z4�?,             O@������������������������       ��5��?             ;@������������������������       �4�2%ޑ�?            �A@[       ^                    �?�������?�           X�@\       ]                     �?P����?�           H�@������������������������       ���|�r�?�             w@������������������������       � �e�?�            �q@_       b                    �?@��!�Q�?P           h�@`       a                     �? �ׁsF�?            y@������������������������       ����C-��?�            �n@������������������������       ���X8��?^            @c@c       d                     �? >��@�?M            @_@������������������������       �        +            @Q@������������������������       ��h����?"             L@f       q                     �?t�G����?�           ��@g       n                    �?кM��K�?�           p�@h       k                    �?�6?JS�?M           �@i       j                    �?��S�ۿ?*            ~@������������������������       �ףp=
�?             $@������������������������       �P&����?%           `}@l       m                    �?H�XA��?#           �}@������������������������       �                     @������������������������       �T�5��%�?            �}@o       p                    �?���?k            �c@������������������������       �                     @������������������������       � ���J��?i            �c@r       y                    �?�>�Y�?�           @�@s       v                    �?�5��JQ�?�           ��@t       u                    �?�LQ�1	�?             7@������������������������       �؇���X�?             ,@������������������������       ������H�?             "@w       x                    �?����$�?|           (�@������������������������       ������?�            0x@������������������������       ��|K��2�?�             p@z       {                    �? 7���B�?B             [@������������������������       �                     @������������������������       ���FM ò?A            @Z@}       �                    �?��iP!�?�           ��@~       �                     �?�	j*D�?�           �@       �                    �?N����?�           H�@�       �                    �?r�q��?             >@������������������������       �P���Q�?             4@�       �                    �?���Q��?             $@������������������������       �      �?              @������������������������       �      �?              @�       �                    �?V�� N��?�           X�@�       �                    �?Z�;nP��?�           p�@������������������������       ��+T{g�?�             w@������������������������       �������?�            �o@������������������������       �L=�m��?(            �N@�       �                    �?x�r���?           �{@�       �                    �?8�Z$���?             *@������������������������       ��<ݚ�?             "@������������������������       �                     @�       �                    �?�fI���?           �z@������������������������       �                     �?�       �                    �?V]�t-��?           �z@�       �                    �?���V��?�            �v@������������������������       ��ǙG=D�?�            @k@������������������������       �Z�/�j��?_            �b@������������������������       �����X�?&            �O@�       �                    �?��C����?�           @�@�       �                     �?��?���?�           ��@�       �                    �?n�C�^��?�            @x@�       �                    �?�r����?             .@������������������������       �                     @������������������������       ��<ݚ�?             "@�       �                    �?Xf�f��?�            Pw@������������������������       ��q���?}             h@������������������������       �������?b            �f@�       �                    �?�.�KQu�?�            �p@�       �                    �?r�����?k            @f@������������������������       �                     @������������������������       ���Uf)�?e            `e@�       �                    �?`Y���?:            �V@������������������������       �                     @������������������������       �v ��?6            �U@�       �                    �?d�� H��?c            �b@������������������������       �        
             ,@�       �                     �?�ZbE���?Y             a@������������������������       �h+�v:�?.             Q@������������������������       ����=�/�?+            @Q@�       �                    �?�r2}�?]           ��@�       �                    �?��g���?;           
�@�       �                    �?�:����?�           ؄@�       �                     �?̌WZ�}�?K            �^@�       �                    �?^������?            �A@������������������������       �      �?             8@������������������������       �                     &@�       �                    �?����!p�?7             V@������������������������       ��U�=���?$            �P@������������������������       �                     6@�       �                     �?|�l�]V�?O            �@�       �                    �?�!�"���?�            �p@�       �                    �?l@!���?{            @i@�       �                    �?Z�K�D��?s            �g@�       �                    �?X��ݥ��?g             e@������������������������       ����la��?J            �\@������������������������       ��+$�jP�?             K@������������������������       �                     3@������������������������       �                     ,@�       �                    �?Z���c��?'            �O@������������������������       ���2(&�?             F@�       �                    �?p�ݯ��?             3@������������������������       ��z�G��?             $@������������������������       �                     "@�       �                    �?�B�R���?�            pq@�       �                    �?~���L0�?�            �n@�       �                    �?X<ev5�?z             h@�       �                    �?:v�S��?s            �f@������������������������       �V������?_            �b@������������������������       ����Q��?            �A@������������������������       �                     $@�       �                    �?���c���?!             J@������������������������       �      �?             H@������������������������       �                     @�       �                    �?�IєX�?             A@������������������������       ��r����?             .@������������������������       �        
             3@�       �                     �?�W�~*t�?�           Ԥ@�       �                    �?tʭ��a�?7           �@������������������������       �                     @�       �                    �?,��M:x�?1           �@�       �                    �?P�� �?�           P�@�       �                    �?����w�?Q           �@������������������������       ������?k            �e@������������������������       �X�V��и?�            @w@������������������������       ����N8�?D            @Z@�       �                    �?� �Gx�?�           ��@�       �                    �?��a�!��?           `x@�       �                    �?@��Cܞ�?�            �t@������������������������       �        A            �X@������������������������       �؞�z�̼?�            @m@������������������������       ��q�q�?,            �L@�       �                    �? ,��-�?�            �m@�       �                    �?�i�y�?v            �g@������������������������       �                    �E@������������������������       ����(-�?[            @b@������������������������       ���[�p�?"            �G@�       �                    �?E�B>��?j           ��@�       �                    �?8ӄ�:�?�           $�@�       �                    �?�醵5��?           ��@������������������������       �                     @�       �                    �?���oǾ?           ȉ@�       �                    �?���\�C�?o           ȁ@������������������������       ���<b�ƥ?w             g@������������������������       ��s�c���?�            x@�       �                    �?     ^�?�             p@������������������������       ��i�y�?)            �O@������������������������       � E59|�?w             h@�       �                    �?6��L�?}            `i@������������������������       ���}����?R            �`@������������������������       �^������?+            �Q@�       �                    �?��%�r�?�            �u@�       �                    �?�\�)G�?�            �p@������������������������       �0�,���?'            �P@������������������������       �< 
2��?�            `i@������������������������       ���Q���?0             T@�                          �?tM����?"	           V�@�                            �?�h�k1P�?�           ��@�       �                    �?�^x�0��?m           x�@�       �                    �?p֤���?�            �u@�       �                    �?�t����?�            �m@������������������������       �����#��?�             i@������������������������       ����@��?            �B@������������������������       � '��h�?E            @[@�       �                    �?`O����?�            �n@������������������������       �5�wAd�?T            �`@������������������������       �        9            �[@                         �?��R[s�?�           h�@                         �?\�����?�           �@                         �?f�{�S �?�           ��@������������������������       ��$d�ď�?*           �}@������������������������       �Բ r��?^             c@                         �?��S���?,            �R@������������������������       ��KM�]�?             C@������������������������       ��?�|�?            �B@	      
                   �?���G��?�            �u@������������������������       �8Fi#]�?�            �q@������������������������       �(;L]n�?+             N@      !                   �?.;[����?(           ��@                         �?B0�8���?p            �e@                         �?�2����?$            �K@                          �?      �?             8@������������������������       ��C��2(�?             &@������������������������       ��n_Y�K�?             *@                          �?��a�n`�?             ?@������������������������       �ףp=
�?             $@                         �?�����?             5@������������������������       ��8��8��?             (@������������������������       ������H�?             "@                         �?P���Q�?L             ^@                         �?x�}b~|�?&            �L@                          �?dP-���?            �G@������������������������       �@4և���?             ,@������������������������       ��C��2(�?            �@@                          �?ףp=
�?             $@������������������������       �                     @������������������������       �r�q��?             @                           �? ������?&            �O@������������������������       �                     <@������������������������       ���?^�k�?            �A@"      -                   �?��V]O�?�           L�@#      &                   �?���W"��?E           �@$      %                    �?�f��>�?�           H�@������������������������       ��J�ۈ�?�            `q@������������������������       �h!�'nf�?�            0u@'      *                   �?L�[2[
�?�           ��@(      )                    �?���g<�?�            �q@������������������������       � 	��p�?Z             b@������������������������       ��#-���?X            �a@+      ,                    �?�<�� �?           �{@������������������������       �L�[2[
�?r            �f@������������������������       �T��o��?�            Pp@.      5                   �?0��Nhk�?s           ��@/      2                   �?���w��?�            Py@0      1                    �?X�<ݚ�?�            �r@������������������������       �� �	��?X            @_@������������������������       ����EH��?j            �e@3      4                    �?�>���?<             [@������������������������       ��û��|�?             G@������������������������       ��g�y��?!             O@6      7                    �?p�EG/��?u            �g@������������������������       ���.���?5            �U@������������������������       �������?@            �Y@9      �                    �?��Y�?�+           &�@:      W                   �?D���O�?�           q�@;      F                   �?Ȱl�?1	           4�@<      A                   �?�A�$�ʚ?�           ��@=      @                   �? ��s`�?�            r@>      ?                   �?@�j;��?Y            �a@������������������������       �                     @������������������������       ����}<S�?W            @a@������������������������       �        T            `b@B      E                   �?�='�1Nu?�           ��@C      D                   �?�i�%��?�            `i@������������������������       �                     2@������������������������       � S5W�?|             g@������������������������       � �^��l?_           ��@G      P                   �?p�"�0�?�           ��@H      K                   �?R��MG��?�           L�@I      J                   �?�hO�B�?�            ps@������������������������       ��6�`g�?g            �e@������������������������       ��!���?R             a@L      M                   �?ȸ�{J^�?�           ��@������������������������       � ��fί�?�            `y@N      O                   �?�"%�a�?�            `x@������������������������       �                     �?������������������������       �0�]]#�?�            Px@Q      T                   �?�i�T�?�           ��@R      S                   �?�4}5�?�             r@������������������������       ���[�A�?Q            �^@������������������������       �d}h���?i             e@U      V                   �?����?8           �@������������������������       �8��cV�?,           �|@������������������������       �Xe�&��?           ��@X      m                   �?ԙ@s��?c	           ��@Y      f                   �?`+*���?t           ��@Z      _                   �?z�G�z�?C           @@[      ^                   �?�� �JH�?�            �m@\      ]                   �?�|���?5             V@������������������������       �                    �H@������������������������       � ���J��?            �C@������������������������       �        `            �b@`      c                   �?      �?�            �p@a      b                   �?�{ /h��?j            �c@������������������������       �ҳ�wY;�?;            @U@������������������������       �:%�[��?/            �Q@d      e                   �?f<t=9%�?D             [@������������������������       ��̚��?'            �N@������������������������       �z�J��?            �G@g      j                   �?�e"���?1           Ћ@h      i                   �?��!����?           �y@������������������������       �X��Oԣ�?�             o@������������������������       �@�#����?e             d@k      l                   �?@[���?)           ~@������������������������       �$�q-�?�            @p@������������������������       ���Au5a�?�            �k@n      y                   �?������?�           Ң@o      t                   �?���PXY�?�           ȃ@p      s                   �?fP*L��?�            �p@q      r                   �?�+e�X�?,            �R@������������������������       �:	��ʵ�?            �F@������������������������       ��q�q�?             >@������������������������       ��? Da�?j            �g@u      x                   �?,���i�?�            w@v      w                   �?�z<�L�?^            `b@������������������������       �        4            �T@������������������������       �D������?*            @P@������������������������       ��g+��@�?�            �k@z                         �?���l��?o           ��@{      ~                   �?�Ŗ�Pw�?f           @�@|      }                   �?�Ru߬Α?L            �\@������������������������       �                     @������������������������       ���wڝ�?H            @[@������������������������       ��1���܋?           `{@�      �                   �?P����N�?	            �@�      �                   �?��]�ӵ�?�            �t@������������������������       �                      @�      �                   �?�_�ܹ��?�            �t@������������������������       �      �?1             R@������������������������       ��^龆��?�             p@�      �                   �?��v����?#           ��@������������������������       �T�iA�?P            �a@������������������������       ������t�?�           ��@�      �                   �? ���N�?          ���@�      �                   �?t�e��P�?F           �@�      �                   �?$>:1���?�           z�@�      �                   �?�w�\Q�?�           (�@�      �                   �?�����?            `|@������������������������       �        )             O@�      �                   �?0��X�t�?�            �x@������������������������       �Xc!J�ƴ?E            �]@������������������������       ��(�T[X�?�             q@�      �                   �?H�㸪�?}           �@�      �                   �?d-�Q�?�            pq@������������������������       ��U�!��??            @X@������������������������       �t]����?m            �f@�      �                   �?HQ�k�?�           h�@�      �                   �?��ف�"�?�            �r@������������������������       �                     �?������������������������       �D��F�5�?�            �r@�      �                   �?�����η?            |@������������������������       �                     @������������������������       ��6�4��?           �{@�      �                   �?b�=#O�?!           `�@�      �                   �?�4�'�@�?            ��@������������������������       ��\����?f            `d@������������������������       � ��[��m?�           �@�      �                   �?8௷�c�?           $�@�      �                   �?�z/sT�?�            @v@������������������������       �0B��D�?G            �]@������������������������       �z�����?�            �m@�      �                   �?��q㹤�?           ��@������������������������       ��X�<ݺ?            {@������������������������       �8�'�h׷?           Ԓ@�      �                   �?V�����?�           D�@�      �                   �?���4��?k            �@�      �                   �?��wڝ�?A            @[@������������������������       �                     �?�      �                   �?`�߻�ɒ?@             [@������������������������       ��Ń��̧?             E@������������������������       �        %            �P@�      �                   �?B2�'5��?*           p}@������������������������       �                     �?�      �                   �?��G�߈�?)           `}@�      �                   �?�&z�,�?Q            @^@������������������������       ��q�q�?,            �O@������������������������       ��c�Α�?%             M@�      �                   �?����e��?�            �u@������������������������       ������H�?t            �g@������������������������       �ףp=��?d             d@�      �                   �? 
��р�?           h�@�      �                   �? ��]���?�            �p@�      �                   �?v���a�?4            @R@������������������������       �                     ?@������������������������       �0,Tg��?             E@�      �                   �?��D���?w             h@������������������������       �        X             c@������������������������       ��G�z��?             D@�      �                   �? E59|�?r           �@������������������������       ��1Y�I��?�            �l@������������������������       ���K�Φ?�            �u@�      �                   �?,A����?�	           8�@�      �                   �?`�j���?Q           ��@�      �                   �? ���g=�?�            �i@�      �                   �?&[i`��?3            �U@������������������������       � �h�7W�?            �J@������������������������       ���.k���?             A@������������������������       � �q�q�?T             ^@�      �                   �?@����?�            �@�      �                   �?`�LVXz�?�            �h@������������������������       �                     <@������������������������       �`��>�ϗ?q            @e@�      �                   �?\G2��?G           �@������������������������       ���7Y��?D            �[@�      �                   �?���@�ϻ?           �x@������������������������       �                     @������������������������       �@��S�$�?�            �x@�      �                   �?H2rY��?o           �@�      �                   �?@�Dw�@�?�           t�@������������������������       � ����?+            @P@������������������������       � "���?�           p�@�      �                   �?@��Y��?�           ��@�      �                   �?�� d,l�?�            `v@������������������������       ��	j*D�?             J@������������������������       ��X�<ݺ?�             s@�      �                   �?x�;����?�           �@������������������������       ���8AK�?}            �g@������������������������       �@(8�?B           �@q�tq�bh�h"h#K �q�h%�q�Rq�(KM�KK�q�hQ�B�      �i�@    @��@    ���@     ��@    ���@     �@     �|@     �}@     @|@     �}@     �w@     `t@     @l@      l@     �b@     @Y@      S@     @b@      @      �?       @              @      �?       @               @      �?    ���@     ��@    �e�@     (�@    �@�@     �t@     ��@      `@     ��@     @^@     �@     �U@     ��@     �B@     �W@      �?     @T@      �?      ,@             ��@      B@     �@      =@     @q@      @      u@      I@      m@     �F@      ?@      "@     @i@      B@     �Y@      @      @              Y@      @     �K@      A@      D@      *@               @      D@      &@      .@      5@     @[@      @     �C@      @      9@      @      @              6@      @      ,@      @      �?              *@      @     �Q@            ���@     @i@     �@     @Y@     �`@             m�@     @Y@     T�@      @     ��@      @     ��@             ��@     �W@     X�@     �R@     ��@      B@     ��@      C@     pq@      4@     L�@     @Y@     ԓ@      @     �@      @      7@             0�@      @     ��@      �?      4@              �@      �?     ~@      �?     �X@             Ę@     �W@      "@             ��@     �W@     �@     �S@     x�@      E@     P�@     �B@     �e@      .@     ��@     �s@     ԕ@     �e@     �m@     �c@     �k@     @\@     �a@      U@     �[@      @@     �@@      J@     @S@      =@      M@      0@      3@      *@      3@     �E@      &@      0@       @      ;@     �@      0@     ��@      &@     �v@      @     0q@      @     @�@      @     �x@      @     �n@      �?     �b@      @      _@      �?     @Q@             �K@      �?     T�@     �a@     `�@      Q@     �@      P@      |@      @@      "@      �?     p{@      ?@     �{@      @@      @             �{@      @@     `c@      @      @              c@      @     �@     �R@     ��@     �Q@      4@      @      (@       @       @      �?     �@      Q@     �u@      E@      m@      :@      Z@      @      @             @Y@      @     �@     H�@     �@     @v@      ~@     �l@      @      9@      �?      3@      @      @      @      @      �?      �?     �}@     �i@     �z@     `h@     �p@     @Y@     �c@     �W@      I@      &@     �s@     @_@       @      &@       @      @              @     �s@     �\@      �?             �s@     �\@     �p@      X@     �c@     �M@      \@     �B@     �F@      2@     0z@     Px@     u@      t@      g@     `i@       @      *@              @       @      @     �f@     �g@      W@      Y@     �V@     �V@      c@     @]@     �Z@      R@              @     �Z@     @P@      G@     �F@              @      G@      D@     �T@     @Q@              ,@     �T@     �K@      E@      :@      D@      =@     n�@     ��@     z�@     @�@     `l@     �{@      1@     �Z@      (@      7@      (@      (@              &@      @     �T@      @     �N@              6@     @j@     �t@     �`@     �`@      ^@     �T@      ^@      Q@     @Y@      Q@     �L@      M@      F@      $@      3@                      ,@      *@      I@      @      C@      @      (@      @      @              "@     @S@     @i@     �R@     @e@      Q@     @_@      M@     @_@      F@      Z@      ,@      5@      $@              @     �F@      @     �F@      @               @      @@       @      *@              3@     ��@      q@     ��@     �W@      @             x�@     �W@     �@     �F@     h�@      4@     �e@      �?     v@      3@      T@      9@     �@     �H@     Pv@     �@@     �s@      ,@     �X@             �k@      ,@      C@      3@     �k@      0@     �f@      @     �E@             �a@      @     �B@      $@     Ԓ@     @f@     `�@     @_@     H�@     �J@      @              �@     �J@     h�@      F@     �f@      @     �u@      D@     �n@      "@     �N@       @     @g@      @     ``@      R@     @U@      H@      G@      8@     �r@     �J@     �n@      :@     @P@       @     `f@      8@     �J@      ;@     b�@     �@     ��@     ,�@      q@     �s@     �@@     �s@      <@     @j@      4@     �f@       @      =@      @      Z@     �m@      @      `@      @     �[@             �p@     `�@     �h@     �@     �c@     �}@      1@     �|@     �a@      &@      D@     �A@      @      A@      B@      �?     �Q@     q@      *@     �p@      M@       @     L�@     x�@      J@     �^@      G@      "@      2@      @      $@      �?       @      @      <@      @      "@      �?      3@       @      &@      �?       @      �?      @     �\@      @      J@      @     �E@      �?      *@      @      >@      �?      "@              @      �?      @      �?      O@              <@      �?      A@     |�@     @{@     8�@     `f@     0�@     �X@     �m@      D@     �q@     �M@     @�@      T@     pp@      6@     �`@      $@      `@      (@     x@      M@     @d@      4@     �k@      C@     u@     p@     �k@     �f@     �d@     �`@     �Q@     �K@     �W@     @S@      M@      I@      <@      2@      >@      @@     �\@     �R@     �L@      =@     �L@      G@     ��@     \�@     ��@     ��@      u@     ��@      ,@     H�@      (@     Pq@      (@     @`@              @      (@     �_@             `b@       @     �@      �?     @i@              2@      �?      g@      �?     ��@     @t@     l�@     `g@     ��@     �[@      i@     �P@     @[@      F@      W@     @S@     x�@      B@      w@     �D@     �u@              �?     �D@     �u@      a@     x�@     @Q@     �k@     �@@     @V@      B@     �`@      Q@     �@      1@     �{@     �I@     H�@     Px@     ��@     �e@      �@      Y@      y@      �?     `m@      �?     �U@             �H@      �?      C@             �b@     �X@     �d@      M@     �X@      >@     �K@      <@     �E@     �D@     �P@      2@     �E@      7@      8@     �R@     ��@      D@     w@      <@     �k@      (@     �b@      A@     �{@      4@      n@      ,@     �i@     �j@     $�@     �U@     �@      E@     �k@      2@     �L@       @     �B@      $@      4@      8@     �d@     �F@     @t@      ?@      ]@             �T@      ?@      A@      ,@      j@      `@     ��@      @      �@      �?     @\@              @      �?      [@      @     0{@      _@     0�@     �D@     0r@               @     �D@     r@      2@      K@      7@     `m@     �T@     H�@      M@     �T@      9@     ��@     H�@     �@     �@     �@     �w@      �@     �f@     X�@      $@     �{@              O@      $@     �w@      @     @\@      @     �p@     @e@     Њ@     �\@     �d@     �H@      H@     �P@      ]@     �K@     ��@     �@@     �p@              �?     �@@     �p@      6@     �z@              @      6@     pz@     �h@     ԧ@      @     ��@      @      d@       @     �@      h@      �@     �[@     �n@      >@      V@      T@     �c@     �T@     H�@      8@     �y@     �M@     �@      `@     D�@     �S@     `@      �?      [@              �?      �?     �Z@      �?     �D@             �P@     @S@     �x@              �?     @S@     �x@     �B@      U@      5@      E@      0@      E@      D@     Ps@      5@      e@      3@     �a@      I@     ؈@      =@     �m@      &@      O@              ?@      &@      ?@      2@     �e@              c@      2@      6@      5@     p�@      *@     �j@       @     pu@     �p@     �@     �W@     ��@      8@     �f@      3@      Q@      @      I@      0@      2@      @     �\@     �Q@     �@       @     �h@              <@       @      e@     @Q@     �{@      G@     @P@      7@     �w@              @      7@     0w@      f@     ��@      @     `�@      �?      P@      @     `�@     `e@     �@     �@@     Pt@      0@      B@      1@     r@     @a@     �@     �O@      `@     �R@     �@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       qԆq�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheM�hfh"h#K �q�h%�q�Rq�(KM��q�hm�B�g         F                   �?�����?�e           �@       �                    �?�dƉq��?�D          �D�@       `                    �?`d�y��?:(           ��@                           �?�$p�Z�?K          �O�@       
                    �?��}*_��?G           ��@       	                     �?
��p���?f           ��@                            �?ʽ�C�?�           ��@������������������������       ���͵���?           Pz@������������������������       ��L�lRT�?�            �p@������������������������       �X������?�            �p@                           �?�������?�            �v@                           �?\����?�            �u@                           �?,d��?�            �t@                           �?0�`G�r�?�            `t@                            �?�.(�i��?Y            �b@                           �?P�Lt�<�?B            �\@������������������������       ��|1)�?;            �Z@������������������������       �                      @                           �?��G���?            �B@������������������������       ��'�`d�?            �@@������������������������       �                     @������������������������       �        p            �e@                           �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             ,@������������������������       �                     4@       K                    �?����Q�?           ��@       <                    �?�5)0g�?�          ���@       /                    �?�o�P���?�          �W�@       &                     �?�Τ�F�?�           q�@        #                    �?`��f�?�           f�@!       "                    �?X��8�y�?           (�@������������������������       �le}����?l           �@������������������������       �z�G�z�?            �A@$       %                    �?��ŽR��?)           ��@������������������������       � ��f�r?W           ,�@������������������������       �H�joѸ?�           �@'       ,                    �?X�g>���?�           ��@(       )                    �?w\e1��?#           H�@������������������������       �                     �?*       +                    �?��4��?"           @�@������������������������       ��uD����?�             m@������������������������       �@[�Ik��?�           ��@-       .                    �?0ia�2ͬ?�           ��@������������������������       ��}�+r��?             3@������������������������       �Bli�/�?�           �@0       7                    �?��F�D�?1
           >�@1       4                    �?����SS�?
           ,�@2       3                     �?h(I�1ɶ?           py@������������������������       ���ݶ3�?�            r@������������������������       ��j��b�?K            �]@5       6                     �? D,�T?�           И@������������������������       �        �           L�@������������������������       � P�@��p?3           ~@8       9                    �?R�_�f�?'           �@������������������������       �                    �E@:       ;                     �?�Q����?           ��@������������������������       ��DC'j�?c           p�@������������������������       ������?�           `�@=       D                    �?�B!Ae�?�           ��@>       A                     �? �&�eZ�?�             s@?       @                    �?蹱f
@�?z            �e@������������������������       ��iyw	
�?\            �`@������������������������       �                    �C@B       C                    �?0�!F��?T            �`@������������������������       ���F�D�?;            �X@������������������������       �l��\��?             A@E       H                     �?6Pc���?           �{@F       G                    �?�vc%��?�            Pp@������������������������       ��`⯛��?e            �c@������������������������       �<=�,S��?@            @Z@I       J                    �?�N��M��?n             g@������������������������       ��n_Y�K�?H            @]@������������������������       �.Lj���?&             Q@L       W                    �?�B��el�?i           ��@M       T                    �?�&�5y�?            {@N       Q                    �?x�}b~|�?�            `u@O       P                     �?�w�r��?2            @S@������������������������       ���s����?             E@������������������������       ���
P��?            �A@R       S                     �? ���Sr�?�            �p@������������������������       �        f             e@������������������������       ���8�$>�?9            @X@U       V                     �?hl �&�?5             W@������������������������       �`'�J�?            �I@������������������������       ���Y��]�?            �D@X       ]                    �?$��t�r�?c           �@Y       Z                    �?%Xhqv�?5           �}@������������������������       �                     &@[       \                     �?@��z��?.           @}@������������������������       � �(�V�?�            �p@������������������������       ������?}            �h@^       _                     �?�v:���?.             Q@������������������������       �^������?            �A@������������������������       �����e��?            �@@a       �                    �?�$ �?�
           E�@b       �                    �?��9[��?`           $�@c       r                    �?��5V�?�           ��@d       o                    �?z�G�z�?^            `c@e       j                     �?�e+��?K            @^@f       i                    �?��
ц��?            �C@g       h                    �?����"�?             =@������������������������       �`�Q��?             9@������������������������       �      �?             @������������������������       �                     $@k       n                    �?ĴF���?0            �T@l       m                    �? wVX(6�?/            @T@������������������������       ���(\���?.             T@������������������������       �                     �?������������������������       �                     �?p       q                     �?l��\��?             A@������������������������       �                     "@������������������������       �H%u��?             9@s       ~                    �?K��J>�?�           P�@t       {                    �?DX�\��?           �z@u       x                     �?\������?�             t@v       w                    �?E����?\            `b@������������������������       ��/���??            �Y@������������������������       ��������?             F@y       z                    �?��M$i�?p            �e@������������������������       ��>z���?W             a@������������������������       ���
ц��?            �C@|       }                     �?�ջ����??             Z@������������������������       ���hJ,�?             A@������������������������       �b�h�d.�?'            �Q@       �                    �? �z�[�?�           P�@�       �                    �?�O4R���?I           ��@�       �                     �?�s��;�?�            @v@������������������������       �@�Gpm��?p             g@������������������������       ������?k            `e@�       �                     �?�B:�g�?n            �e@������������������������       �        @             [@������������������������       �����e��?.            �P@�       �                     �?�zvܰ?7             V@������������������������       �                    �B@������������������������       ��IєX�?            �I@�       �                     �? p}U�?w           �@�       �                    �?�c�ZB�?�             y@�       �                    �?�_%����?�            �l@������������������������       �                     8@������������������������       � �O���?~            �i@�       �                    �?`<�Gf�?o             e@������������������������       �                     "@�       �                    �?      �?i             d@������������������������       �`Ӹ����?             �F@������������������������       ���x$�?I            �\@�       �                    �?�\�2�q{?|           ��@�       �                    �?@Fd�4�?�            �u@������������������������       �        $            �K@������������������������       � I!�}�?�            �r@������������������������       �        �            �n@�       �                    �?>�ÌG�?�           f�@������������������������       �                      @�       �                     �?�[�#K�?�           b�@�       �                    �?�z�6�?�           x�@�       �                    �?�#�S�`�?�           ��@�       �                    �?���}<S�?             7@������������������������       �                     3@������������������������       �      �?             @�       �                    �?�P�D�߷?�           8�@�       �                    �?�NWm��?�           (�@������������������������       ��q�q�?�             x@������������������������       ��J��?�            �l@������������������������       �@3����?i            @d@�       �                    �?    ���?�             p@�       �                    �?^n����?u            �f@������������������������       ��j�8���?P            �\@������������������������       ��y(dD�?%            @P@������������������������       ��I�w�"�?.             S@�       �                    �?��<^�?�           L�@�       �                    �?zL��#��?(           H�@�       �                    �?�u�[A��?�           8�@�       �                    �?����?           0{@������������������������       �                      @������������������������       �85�}C�?           �z@�       �                    �?�|1)��?�            �j@������������������������       �                      @������������������������       ��IJ��?�            @j@�       �                    �?f�Ý��?�            @l@������������������������       �П[;U��?t            �e@������������������������       ���WV��?"             J@�       �                    �?�7�r��?�            �r@�       �                    �?\� ���?�            �h@������������������������       �                      @������������������������       ���`ۻ��?�            �g@������������������������       ���.k���?=            �Y@�                          �?V���v��?�           ��@�       �                    �?V�p����?�           ��@�       �                    �?ڨ�Nޯ�?!	           �@�       �                    �?l�a+\5�?O           $�@������������������������       �                     @�       �                    �?�k��f��?M           �@�       �                    �?�������?�            �w@�       �                     �?�[�|Tc�?�            �o@�       �                    �?�('+��?]            �a@������������������������       ����c�?W            �`@������������������������       ��z�G��?             $@�       �                    �?p�s(���??            �[@������������������������       ��	��)��?:            �Y@������������������������       �؇���X�?             @�       �                     �?R�c���?S             `@�       �                    �?*c̕6�?9            �U@������������������������       �j(���?4            @S@������������������������       �ףp=
�?             $@�       �                    �?����X�?             E@������������������������       �<ݚ)�?             B@������������������������       �r�q��?             @�       �                    �?��3EaǼ?^            �@�       �                    �?�_�V��?�           �@�       �                     �?���;���?�           h�@������������������������       ����.�*�?�            �u@������������������������       � ��(�?�            0q@�       �                     �?�:�^���?           ��@������������������������       ��n;I�"�??           0@������������������������       ��+I�9��?�            @v@�       �                     �?�2�~w�?�           0�@�       �                    �?H�*�ɺ?�           ��@������������������������       � ��7��?�            �n@������������������������       �D�0(?c�?           �z@�       �                    �?��Wv��?            {@������������������������       �        e             c@������������������������       ��5���?�            pq@�       �                    �?��֖�N�?�           ��@�       �                    �?�)f5��?            �y@�       �                     �?pY���D�?�            �s@������������������������       � I!�}�?Z            �b@������������������������       � �q�q�?g             e@�       �                     �?`�q�0ܴ??            �W@������������������������       �@4և���?$             L@������������������������       �                     C@�       �                    �?:"Z��?�            �u@�       �                     �?���j��?�            �l@������������������������       ��%o��?N            �`@������������������������       ��q�Q�?@             X@�       �                     �?�����?D            �\@������������������������       �v�_���?.            �S@������������������������       ���R[s�?            �A@�                          �?"��5��?�
           ,�@�       �                     �?�9Y�\�?�           �@�       �                    �?�Ba[L�?]           ��@�       �                    �?�CR��?�            �@�       �                    �?b�X�O��?�            @u@������������������������       �0�ڂcv�?�            `j@������������������������       �0Ƭ!sĮ?V             `@�       �                    �?4�R�f�?�             s@������������������������       ����!pc�?             &@������������������������       �L��n��?�            Pr@�       �                    �? @|���?�           ��@������������������������       �        O           @�@������������������������       ��������?r            �f@�                          �?�_|0�?x           P�@�                           �?���b���?�           Ԙ@�       �                    �?"��ք�?\           ��@������������������������       �h�����?           @z@������������������������       �(;L]n�?N             ^@������������������������       ��K�-l\w?�           d�@                         �?a�^4�?�           ��@                         �?�o��gn�?�            �t@������������������������       �����X�?             @������������������������       �P6=���?�            Pt@������������������������       �>��8z��?�            pr@                          �?�(���?�            �@                         �?0lؕ���?�            �w@	                         �?>A�F<�?�            �l@
                         �?v�X��?             F@������������������������       ����y4F�?             C@������������������������       �r�q��?             @                         �?��3EaǼ?v             g@������������������������       �                    �D@������������������������       �$�q-�?[            �a@                         �?��F��?^            `c@������������������������       �        F            �\@������������������������       �� ��1�?            �D@                         �?:�=�a��?           Pz@                         �?�8�So��?�            @n@                         �?$��m��?3            �S@������������������������       ������?             C@������������������������       ��(\����?             D@                         �?����?a            �d@������������������������       �      �?             @������������������������       � �\���?]            �c@                         �?d��ϸ�?t            `f@������������������������       �`o��b�?S             _@������������������������       �<|ۤ$�?!            �K@      5                   �?��z���?�           ��@      *                   �?�����?�           ޡ@       %                    �?<����?�            pu@!      $                   �?,�[I'��?u            �g@"      #                   �?t�F�}�?=            �Y@������������������������       �#z�i��?            �D@������������������������       ���v$���?&            �N@������������������������       �        8            �U@&      )                   �?���u��?]            `c@'      (                   �?~���L0�?;            �X@������������������������       �����X�?             E@������������������������       �        $             L@������������������������       �0�)AU��?"            �L@+      2                   �?��Wv��?�           `�@,      /                   �?,����?2           p}@-      .                    �? �ղ?�            �v@������������������������       �ȑ����?H            @]@������������������������       ��,_���?�             o@0      1                    �?@��!�Q�?B            @Z@������������������������       �                     H@������������������������       �0�)AU��?&            �L@3      4                    �?@B����?�           �@������������������������       �                   `{@������������������������       ���Ij�?�           ,�@6      ?                   �?���o^��?           <�@7      8                   �?4Qi0���?�           �@������������������������       �        	             *@9      <                   �?�[Y��.�?�           ��@:      ;                    �?�%IM��?�            �q@������������������������       �(32v�c�?q            `d@������������������������       �H��ԛ�?N            �]@=      >                    �?t��x��?           �{@������������������������       ���I�� �?q            `f@������������������������       ����L:�?�            �p@@      C                    �?��f|��?'           �z@A      B                   �?F��{�?~            �g@������������������������       �^l��[B�?$             M@������������������������       ��c��{-�?Z            ``@D      E                   �?^n����?�             n@������������������������       ��d�����?"            �L@������������������������       ��q�q�?�            �f@G      �                   �?���ž�?�            ��@H      �                   �?��āι�?�           S�@I      f                   �?�,X����?8           L�@J      W                   �?���K���?            0�@K      R                    �?���C��?#            �J@L      O                   �?��� ��?             ?@M      N                   �?$�q-�?
             *@������������������������       �                     "@������������������������       �      �?             @P      Q                   �?r�q��?             2@������������������������       �                     $@������������������������       �      �?              @S      V                   �?�C��2(�?             6@T      U                   �?�q�q�?             @������������������������       ��q�q�?             @������������������������       �                     @������������������������       �        	             0@X      _                   �?B�,rVL�?�           \�@Y      \                   �?��}V�?+           ��@Z      [                    �?�P�p��?[           ��@������������������������       ��H�7��?�            pu@������������������������       ��<ݚ�?�            �g@]      ^                    �?��}*_��?�            @t@������������������������       ��Q�N��?r            �f@������������������������       ����|���?^            �a@`      c                    �?�T��?�           ��@a      b                   �?{I��%�?           �{@������������������������       ��������?�            Pq@������������������������       �d�m�v��?d            @e@d      e                   �?    ��?�             p@������������������������       �����X�?j            �e@������������������������       �|��?���?7            @T@g      v                   �?�'wݥ�?8           Њ@h      o                   �?�+�$f��??            �X@i      l                    �?X�EQ]N�?            �E@j      k                   �?؇���X�?             5@������������������������       �     ��?	             0@������������������������       �                     @m      n                   �?�C��2(�?             6@������������������������       ��KM�]�?
             3@������������������������       �                     @p      s                   �?lGts��?&            �K@q      r                    �?X�EQ]N�?            �E@������������������������       �@�0�!��?	             1@������������������������       �$�q-�?             :@t      u                    �?�8��8��?             (@������������������������       �                     @������������������������       ������H�?             "@w      ~                   �?��f�-y�?�           ��@x      {                   �?�T��5m�?            y@y      z                    �?�ˍ_��?�            �p@������������������������       �8�A�0��?H            �[@������������������������       �l�a���?_            `c@|      }                    �?�Eǎ\�?\             a@������������������������       ��q�q�?4            �R@������������������������       �`՟�G��?(             O@      �                   �?dT�Z*S�?�            `v@�      �                    �?�Pf����?�            �q@������������������������       ��n\�GZ�?P            �]@������������������������       ���w�T�?q            �d@�      �                    �?�;�vv��?5            @R@������������������������       �      �?             8@������������������������       ��`���?"            �H@�      �                   �?�ܵ�|@�?�            �@�      �                   �?x���s(�?_           �@�      �                   �?T~bl]i�?�           �@�      �                    �?Ddq���?�           p�@������������������������       ��ڊ�e��?�             y@�      �                   �?��2(&�?�            �q@������������������������       �                     �?������������������������       �\�ih�<�?�            �q@�      �                    �?�:�]��?           �|@������������������������       �|�db���?�            �p@������������������������       ��V���?r            �g@�      �                   �?�FVQ&�?�           ,�@�      �                    �?��{V��?V           ��@������������������������       ��g�.�?A           �@������������������������       ���Ujѡ�?           @{@�      �                    �?�|����?1           `}@������������������������       ����}<S�?�            �o@������������������������       �|H�=|k�?�             k@�      �                   �?��wV��?V	           ��@�      �                    �?�d!����?�           ,�@�      �                   �?6����?r           0�@�      �                   �?�����?           pz@������������������������       �                     �?������������������������       ���P����?           `z@������������������������       �D���D|�?m            �c@�      �                   �?P�p�(+�?�           (�@������������������������       �                     @�      �                   �?p���p�?�           ��@������������������������       � >�=���?           `|@������������������������       �pb����?k             g@�      �                    �?8�9�e�?[           b�@�      �                   �?��?�/�?�            �@������������������������       ���D����?�           ��@������������������������       �Dw�&��?�            �j@�      �                   �?��L�?�           ��@������������������������       �P�~(w}�?�           T�@������������������������       �xX7�Ӳ?�            @u@�      �                   �?��QY�q�?�
           0�@�      �                   �?x4�	��?�           І@�      �                   �?��4"�?�?�            pr@�      �                    �?�[�}r�?Z            ``@�      �                   �?*O���?/             R@������������������������       �      �?             @������������������������       �.Lj���?,             Q@�      �                   �?:���W�?+            �M@������������������������       �                     @������������������������       ���X��?(             L@�      �                   �?�{��?c            �d@������������������������       �                     2@�      �                    �?:PZ(8?�?X            @b@������������������������       ��������?(             Q@������������������������       ��n_Y�K�?0            �S@�      �                   �?L�A���?           0{@�      �                   �?�Fǌ��?/            �S@������������������������       �        
             1@�      �                    �?0�z��?�?%             O@������������������������       �                     5@������������������������       ���Y��]�?            �D@�      �                    �?��!h
��?�            @v@�      �                   �?>�6�%�?w            `g@������������������������       ��q�q�?7             U@������������������������       ��ԇ���?@            �Y@�      �                   �?�2����?h             e@������������������������       �<=�,S��?0            �Q@������������������������       �X�<ݚ�?8            �X@�      �                   �?�)�=�?	           ��@�      �                    �?��zx�?�           ��@�      �                   �?�X��D�?�             v@������������������������       �tX�}}��?_            �b@������������������������       �؃��)��?�             i@�      �                   �?�T�Z_�?           p{@�      �                   �?��pBI�?Y            @b@������������������������       �                     �?������������������������       ��=x�?X             b@������������������������       �Ur����?�            Pr@�      �                   �?�a!���?            ~�@�      �                    �?���H`�?�           0�@�      �                   �?�O��/�?�            `q@������������������������       �                      @������������������������       ��θV�?�            @q@�      �                   �?�X�<ݺ?            {@������������������������       �                     @������������������������       �X�޻G�?           �z@�      �                    �?x(�I��?^           �@������������������������       �h�⶞e�?�           ��@������������������������       �����;�?n           ��@q�tq�bh�h"h#K �q�h%�q�Rq�(KM�KK�q�hQ�B�       T�@     ��@    ���@    ���@    �b�@     >�@    �Z�@     ��@     �@     �~@     �~@      }@     0y@      r@     �l@      h@     �e@      X@     �V@      f@     0u@      :@     �s@      :@     �s@      (@     �s@      $@     �a@      $@     �[@      @     �Y@      @       @              >@      @      :@      @      @             �e@              @       @               @      @                      ,@      4@             ��@      �@     +�@     H�@     ��@     0p@     ±@     �e@     ��@     �[@     ��@      H@     Ȁ@     �D@      <@      @      �@      O@      �@      @      �@     �M@     ��@     @P@     �@      F@      �?             ��@      F@     �h@      A@     ��@      $@      �@      5@      2@      �?     p�@      4@     ԯ@      U@     ܞ@      4@     @x@      3@     �q@      @     �Z@      (@     ̘@      �?     L�@              ~@      �?     f�@      P@     �E@             �@      P@     ��@      F@     ��@      4@     @e@     0�@      ,@     @r@      "@     �d@      "@     @_@             �C@      @      `@       @     @X@      @      ?@     �c@      r@      V@     �e@     �H@     �Z@     �C@     �P@      Q@     @]@     �F@      R@      7@     �F@     ��@     �f@     �s@     �]@     �s@      >@     �I@      :@      A@       @      1@      2@     Pp@      @      e@             @W@      @      @     @V@       @     �H@      �?      D@     0~@      P@     �|@      5@      &@             �{@      5@     pp@       @      g@      *@      9@     �E@      (@      7@      *@      4@      �@     Ԝ@     ��@     ��@     P�@     Px@      ?@      _@      <@     @W@      5@      2@      &@      2@       @      1@      @      �?      $@              @     �R@      @     �R@      @     �R@      �?                      �?      @      ?@              "@      @      6@     X�@     �p@     �e@     �o@     �c@     �d@     @V@      M@      K@     �H@     �A@      "@      Q@     �Z@     �G@     @V@      5@      2@      1@     �U@      @      =@      (@      M@     �@      *@     @�@      $@     �u@      "@     �f@      @     �d@      @     �e@      �?      [@             @P@      �?     @U@      @     �B@              H@      @       @     ؎@      @     �x@      �?     �l@              8@      �?     �i@      @     �d@              "@      @     `c@       @     �E@      @      \@       @     ��@       @     �u@             �K@       @     `r@             �n@     x�@     P}@       @             p�@     P}@     �@     �k@     ��@      D@      5@       @      3@               @       @     �@      C@     �@     �A@     �v@      3@     �j@      0@     �c@      @     �R@     �f@     �L@     �^@      A@     @T@      7@      E@      2@      M@     ،@      o@     ��@     `f@     ��@      K@      y@     �A@       @             �x@     �A@      h@      3@       @             �g@      3@     @Y@     @_@     �S@      X@      7@      =@     �l@     @Q@     �f@      .@       @             �e@      .@      H@      K@     ��@     ��@     m�@     ��@     �@     x�@     �@     �p@              @     �@     �p@     �p@      \@      e@      U@      [@     �A@     @Y@      @@      @      @     �N@     �H@     �K@      H@      @      �?     @Y@      <@     �Q@      0@      O@      .@      "@      �?      >@      (@      9@      &@      @      �?     �@     @c@     ��@     @V@      �@      *@     Pu@      @     �p@       @     X�@      S@     �|@      B@     �s@      D@     ,�@     @P@     ��@     �B@     @n@       @     Px@     �A@     @y@      <@      c@             `o@      <@     @\@     �@      (@     �x@       @     @s@      �?     `b@      @      d@      @     �V@      @      J@              C@     @Y@     `n@     @P@     �d@      E@      W@      7@     @R@      B@     �S@      ;@      J@      "@      :@     ��@     h�@     ��@     l�@     `|@     Ќ@     �y@      m@      a@     `i@      (@     �h@     @_@      @     0q@      =@       @      @     �p@      :@      E@     ��@             @�@      E@     @a@     `�@     p�@     �`@     ��@     ``@     �y@      .@     Py@      ]@      @      @     X�@     `x@     �m@      r@      F@      @       @     �q@      E@     �Y@      h@     `z@     �w@     @h@     �g@     @g@      E@      *@      ?@       @      >@      @      �?     �e@      &@     �D@             �`@      &@       @     `b@             �\@       @     �@@     �l@      h@     �i@      C@     �I@      ;@      (@      :@     �C@      �?      c@      &@      @      @     �b@       @      8@     `c@      �?     �^@      7@      @@     ��@     ��@     �p@     ��@     �a@      i@     �R@     �\@     �R@      <@      ,@      ;@      N@      �?             �U@     @Q@     �U@      Q@      >@      (@      >@      L@              �?      L@     �_@     h�@     �]@     v@      ,@      v@      @     @\@      $@     �m@      Z@      �?      H@              L@      �?       @     �@             `{@       @     �@     ��@     �u@      �@     �P@      *@             ��@     �P@     `p@      4@     �b@      .@     �\@      @     �x@      G@     @d@      1@     `m@      =@      b@     �q@      Q@     @^@      *@     �F@     �K@      S@      S@     �d@      .@      E@     �N@     �^@     £@    ���@     �@     $�@     8�@     ��@     ��@     ��@      @     �G@      @      ;@      �?      (@              "@      �?      @      @      .@              $@      @      @       @      4@       @      @       @      �?              @              0@     p�@     H�@     �@     Pq@     pw@     �c@     �l@     �\@     `b@      E@     �i@      ^@     @\@      Q@     �V@      J@     �z@     @q@     @p@     `g@      f@      Y@     �T@     �U@     �d@     @V@     @_@      I@      E@     �C@     �}@      x@      &@     �U@      @      C@      @      2@      @      *@              @       @      4@       @      1@              @      @     �H@      @      C@      @      ,@       @      8@      �?      &@              @      �?       @     �|@     �r@      p@      b@     �e@     �V@     @P@     �F@     @[@      G@      U@     �J@      I@      9@      A@      <@     �i@      c@      e@     @]@     @R@      G@     �W@     �Q@     �B@      B@      (@      (@      9@      8@     @{@     L�@     �h@     ~�@     �[@     (�@     �R@     �@      B@     �v@     �C@     �n@              �?     �C@     �n@      B@     pz@      3@     @o@      1@     �e@     �U@     Ԕ@      F@     H�@      4@     �~@      8@     �y@      E@     �z@      6@     �l@      4@     �h@     �m@     �@     �V@     ��@     �H@     ��@      C@     x@              �?      C@      x@      &@     �b@      E@     ؂@              @      E@     ��@      4@      {@      6@     `d@     �b@     :�@     �Q@     �@      K@     ؇@      0@     �h@     �S@     l�@     @P@     P�@      *@     pt@     ��@     ��@     �x@     �t@     �f@     @\@      U@     �G@      G@      :@      �?      @     �F@      7@      C@      5@              @      C@      2@     �X@     �P@              2@     �X@      H@      I@      2@      H@      >@      k@     `k@      �?     �S@              1@      �?     �N@              5@      �?      D@     �j@     �a@      ]@     �Q@     �H@     �A@     �P@      B@     �X@     �Q@      F@      :@     �K@      F@      j@     
�@     �F@     P�@      7@     �t@      .@      a@       @      h@      6@     z@      @     �a@              �?      @     �a@      2@     0q@     �d@     6�@      J@     ��@      <@     @o@               @      <@      o@      8@     �y@              @      8@     y@      \@     �@      ?@     ��@     @T@     X�@q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h7Kh8Kh9h"h#K �q�h%�q�Rq�(KK�q�hQ�C              �?q�tq�bhEhUh@C       q�q�Rq�hYKhZh[Kh"h#K �q�h%�q�Rq�(KK�q�h@�C       q�tq�bK�q�Rq�}q�(hKheM�hfh"h#K �r   h%�r  Rr  (KM��r  hm�B�f         F                   �?���=���?|e           �@       �                    �?�0�-$�? E          @O�@       d                    �?�'H��?�(           �@                            �?N�P��?�           Z�@������������������������       ���}��?           0{@                           �?|�ㅚ��?�          ���@       
                     �?��B����?M           @�@       	                    �?���z�?�            Pp@������������������������       �    �S�?�             p@������������������������       �                     @                           �?����V�?�            0p@������������������������       �:u��|2�?�            p@������������������������       �                      @       K                    �?�)�V&�?;          �|�@       "                    �?h^Y�$��?�          ���@                            �?x��;(��?�            v@                           �?����8�?�            �p@                           �?����w�?G            @[@                           �?�&=�w��?F            �Z@                           �?��?^�k�?E            @Z@������������������������       �x�G�z�?9             T@������������������������       �                     9@������������������������       �                     �?������������������������       �                     @������������������������       �        e            �c@                           �?X�EQ]N�?6            �U@                           �?��2(&�?'            �P@                           �?��R[s�?            �A@������������������������       ����!pc�?            �@@������������������������       �                      @������������������������       �                     ?@        !                    �?P���Q�?             4@������������������������       �z�G�z�?             @������������������������       �        
             .@#       :                    �?h ��J��?�           ��@$       /                    �?�v}X@�?�           *�@%       ,                    �?���N��?           H�@&       )                    �?���mas�?�           �@'       (                     �?ۖ�u�?�           �@������������������������       � �-�ظ?`           ��@������������������������       ���:x���?�            �h@*       +                     �?�C�dV�?�            �x@������������������������       ���Z�J�?�            0r@������������������������       ��b�E�V�?>            �Y@-       .                     �?�+e�X�?0            �R@������������������������       �ȵHPS!�?             J@������������������������       �
;&����?             7@0       5                     �?@;'��φ?�	           ��@1       2                    �? �Y�_~?�           ��@������������������������       ��?
i!�?j           H�@3       4                    �? �,?�X?Q           ��@������������������������       �        �           ,�@������������������������       � A��� �?d            @d@6       7                    �? �c���?           d�@������������������������       ��k~X��?�           @�@8       9                    �? �p�?p           ��@������������������������       � ΧZ��?3           0~@������������������������       �����r�?=            �[@;       B                     �?�\��;�?+           ��@<       =                    �?��d*��?+           ��@������������������������       �        &             P@>       ?                    �?Ht��a�?           �@������������������������       �X�aC�U�?�           ��@@       A                    �?�¦�Ư?           X�@������������������������       ���}�?��?c           �@������������������������       �8Fi#]�?�            �q@C       F                    �?hڽD,�?            ��@D       E                    �?=QcG��?            �G@������������������������       �H%u��?             9@������������������������       �                     6@G       H                    �?@�i�q
�?�            �@������������������������       �X�<((�?�           ��@I       J                    �?�ʜ��:�?2           H�@������������������������       ���=��?�           ��@������������������������       �w,�e��?�             k@L       Y                    �?��Y��?h           ��@M       V                    �?�cm)a�?           �{@N       O                    �?�4>�Xb�?�            pv@������������������������       �                     *@P       S                     �?蹱f
@�?�            �u@Q       R                    �?����W�?�            `h@������������������������       ��C��2(�?e            @c@������������������������       �                    �D@T       U                    �?p�`Bh�?c            �b@������������������������       ��r�MȢ?H            �Z@������������������������       ����7�?             F@W       X                     �?ĴF���?2            �T@������������������������       ��S����?             C@������������������������       �`���i��?             F@Z       _                     �?������?I           (�@[       \                    �?*W�C*�?�            �r@������������������������       �z�G�Z�?g             d@]       ^                    �?�7����?]            �a@������������������������       ��ެD��?D            �Y@������������������������       ������?             C@`       c                    �?ޚ)�?�             k@a       b                    �?t]����?p            �f@������������������������       �������?D            �[@������������������������       �"` Y��?,            �Q@������������������������       ��������?             A@e       �                    �?�:l�?�
           T�@f       �                    �?��{-�Z�?           x�@g       x                     �?Q�A+��?�           p�@h       s                    �?n�.P���?�             o@i       l                    �?���k&�?x            �g@j       k                    �?�q�q�?             ;@������������������������       ��	j*D�?             :@������������������������       �                     �?m       p                    �?�cR3?��?g            �d@n       o                    �?
���n<�?H            �\@������������������������       �j%�*R��?;            @W@������������������������       �                     6@q       r                    �? i���t�?            �H@������������������������       ��q��/��?             G@������������������������       �                     @t       w                    �?P̏����?$            �L@u       v                    �?؇���X�?            �H@������������������������       �                     $@������������������������       �:�&���?            �C@������������������������       �      �?              @y       |                    �?��;���?�            `w@z       {                    �? f^8���?B            �Y@������������������������       � ��WV�?2            �S@������������������������       �                     9@}       �                    �?ם�-��?�            �p@~       �                    �?��.k���?y            �i@       �                    �?>(}��?_            �d@������������������������       �b�MKm�?[            `c@������������������������       �                     &@�       �                    �?�s��:��?             C@������������������������       ���
P��?            �A@������������������������       �                     @�       �                    �?��ga�=�?*            �P@������������������������       ��^����?%            �M@������������������������       �                      @�       �                    �?P(_j#��?�           ��@������������������������       �                     $@�       �                     �?`-~���?�           ��@�       �                    �?���O�?�           �@�       �                    �?��z*�o�?�            �s@������������������������       ���<b�ƥ?u             g@������������������������       �        X            �`@�       �                    �?`k�W��?�           H�@�       �                    �?��z	ÿ?           H�@������������������������       �P��B�?�            �w@������������������������       �x�U���?�            �m@������������������������       �      �?i             d@�       �                    �?�DK�%d�?�           ��@�       �                    �?п�#���?8           X�@�       �                    �?p�zٕ`�?�            0r@������������������������       � ���J��?|            `h@������������������������       �      �?6             X@�       �                    �?��SZ��?�           @�@������������������������       �hg� 7��?           �z@������������������������       �$Q�q�?{            �g@�       �                    �?���I�?�            @n@������������������������       ����.�6�?             G@������������������������       ��)���Y�?~            �h@�       �                    �?�Y{~u4�?�           `�@�       �                    �?�:�ǁh�?           ��@�       �                    �? �.��?^           H�@������������������������       �        2            �S@�       �                     �?@=��?,           �}@������������������������       ��M��D`�?�            �h@������������������������       � ��F�}?�            0q@�       �                     �?V>�y	��?�            �r@������������������������       ��"���r�?A            �X@������������������������       �Fx$(�?u             i@�       �                    �?��c��?�            �@������������������������       �                     8@�       �                    �?��p=F�?�           `�@�       �                    �?@���增?�            �x@�       �                     �?p���?C             Y@������������������������       �������?             B@������������������������       �     ��?&             P@�       �                     �?�{Ęd�?�            pr@������������������������       ���x$�?L            �\@������������������������       � Y@��?p            �f@�       �                    �?t�z|�?�            r@�       �                     �?�G�z�?K             ^@������������������������       ��e�,��?&            �M@������������������������       �����5�?%            �N@�       �                     �?�n_Y�K�?l             e@������������������������       ���y�:�?)            �P@������������������������       �Jܤm6�?C            �Y@�                          �?��nh���?�          ���@�       �                    �?��jx+h�?�           �@�       �                    �?��y���?�           J�@�       �                    �? ��h�d�?           ��@�       �                     �? ?,pH!�?t           �@�       �                    �?�@�_
�?           ��@�       �                    �?ox%�:�?�            `k@������������������������       �8����?[            @a@������������������������       �������?0            @T@�       �                    �? *E #�y?�           ȃ@������������������������       � �H~�<x?�            u@������������������������       � �q�	�{?�            �r@�       �                    �?X��Oԣ�?^           p�@�       �                    �?��^@=��?S            ``@������������������������       �      �?              @�       �                    �?�D}1o��?Q             `@������������������������       �`՟�G��?>            @W@������������������������       ��<ݚ�?             B@�       �                    �?@]I��?           �z@������������������������       ��q�q�?�             r@������������������������       �        ^            `a@�       �                    �?�D��z�?�           @�@�       �                    �?��[�Av�?�           ��@�       �                     �?T,��mj�?�           ȅ@������������������������       �<���D�?�            �l@������������������������       �@�R��?$            }@�       �                     �?���N8�?'            �O@������������������������       �>���Rp�?             =@������������������������       �������?             A@�       �                     �?������?�            �u@�       �                    �?�D�e���?k            @e@������������������������       ���x$�?K            �\@������������������������       � �Jj�G�?             �K@�       �                    �?XB���?i            �e@������������������������       ����7�?N            �`@������������������������       �                     E@�       �                     �?�����+�?�           ��@�       �                    �?D�ղ��?�            0p@�       �                    �?v�XԖ�?F            �Z@������������������������       �؀�:M�?            �B@������������������������       ���.N"Ҭ?-            @Q@�       �                    �?*(�"u9�?b             c@������������������������       �io8�?H             ]@������������������������       �                    �B@�       �                    �?v�P��?            }@�       �                    �?X�Cc�?7             U@������������������������       �r�q��?             B@������������������������       �        #             H@�       �                    �?�=A�F�?�            �w@������������������������       �Kb8�į?�            �s@������������������������       � =[y��?)             Q@�       �                    �? ��
̃?�	           ��@�       �                     �?�*�oao�?�           ҡ@�       �                    �? L#Ib?,           ��@������������������������       �        �           ��@�       �                    �? t�)Ї?g            `e@������������������������       �P����?$            �M@������������������������       �        C             \@�       �                    �?������?y           ��@�       �                    �?@PPiP=�?           �@������������������������       ���w#'�?f            `d@������������������������       ��p<L�gw?�           \�@�       �                    �?�|���?q             f@������������������������       �                    �E@������������������������       ����%yU�?T            �`@�       �                    �?�����?�           |�@�       �                     �?`��(�?V            �`@������������������������       �        ,             S@������������������������       ����#�İ?*            �M@�                            �?��Nz�I{?�           `�@������������������������       �                   @|@������������������������       ��Z�H݅�?�           P�@      1                   �?��Qq|�?�
           H�@      "                   �?nK�����?B           ��@                          �?4�exa�?           �@                         �?]]���?U           ��@      	                   �? ��}X�?�           ��@                         �?؇���X�?
             ,@������������������������       ��q�q�?             @������������������������       �                      @
                         �?p�P�2��?�           �@������������������������       ��J��_��?-           �}@������������������������       ��)���Y�?�            `r@                         �?������?i           ��@                         �?�|1)��?           �z@������������������������       �؇���X�?             @������������������������       ��Ñ���?           z@                         �?�L���?Q            �[@������������������������       �                     @������������������������       ��#-���?M            @Z@                         �?���]�?�           |�@                         �?     ��?             @@                         �?"pc�
�?             &@������������������������       �����X�?             @������������������������       �                     @                         �?�G��l��?             5@������������������������       �����X�?             ,@������������������������       �؇���X�?             @                         �?���"���?�           ��@                         �?�R�h��?r           �@������������������������       �(h�M쯿?�            �u@������������������������       �@�p��?�             p@       !                   �?���?x.�?<            ~@������������������������       �R���/�?�            �s@������������������������       �h7�R�
�?f            �d@#      *                   �?�@p��?*           ��@$      '                   �?Tڇ0��?�            �t@%      &                    �?�q�q�?�             k@������������������������       �y�w[��?E            @[@������������������������       ��le����?=            �Z@(      )                    �?��$�4��?G            �]@������������������������       ��1��u�?,            @R@������������������������       ��r����?            �F@+      .                   �?�,��t �?a           (�@,      -                    �?��N`.�?           �{@������������������������       �r٣����?m            �d@������������������������       �x\�Ի�?�            0q@/      0                    �?�u̗C��?F            @[@������������������������       ����j��?             G@������������������������       �b����?'            �O@2      =                   �?� J)IC�?�           8�@3      8                    �?      �?�            �w@4      7                   �?T���O�?�             j@5      6                   �?�KM�]�?h             c@������������������������       �                      @������������������������       �H0sE�d�?f            �b@������������������������       �F�����?'            �L@9      <                   �?r�u���?b            �d@:      ;                   �?ЮN
��?C            @\@������������������������       �                     @������������������������       ��1�`jg�?A            �[@������������������������       �����|e�?             K@>      A                    �?8e�mZ��?�           ��@?      @                   �?��h/���?�            @s@������������������������       ��! �	��?p            �g@������������������������       ��o�Nm��?K            @]@B      E                   �?��q%+�?            z@C      D                   �?H!s��?�            `m@������������������������       �����X�?             @������������������������       ��?�'�@�?�            �l@������������������������       ��o��.�?p            �f@G      �                   �?jYf�?|           ���@H      s                   �?d''!|��?�           ��@I      `                   �?�4|'��?�           ��@J      U                    �?h!�ݒ�?�           x�@K      P                   �?�t����?�           ��@L      M                   �?�C��2(�?             6@������������������������       �                     *@N      O                   �?�<ݚ�?             "@������������������������       �      �?             @������������������������       �z�G�z�?             @Q      T                   �?l`����?�           Ђ@R      S                   �?���{x�?g           ��@������������������������       �
�>Τ�?�            Ps@������������������������       �&��%U�?�             m@������������������������       �r�q��?$             N@V      W                   �?^����?           �z@������������������������       �                     �?X      [                   �?F�E���?           �z@Y      Z                   �?�U�u]�?�            `h@������������������������       ��eP*L��?             &@������������������������       ���wy���?{             g@\      ]                   �?.��$�?�            @m@������������������������       �                     (@^      _                   �?XCwGC�?�            �k@������������������������       ��|G7�?n            �d@������������������������       ��1�`jg�?$            �K@a      h                   �?�Q�Nz2�?           p�@b      g                   �? pƵHP�?             J@c      d                   �?Pa�	�?            �@@������������������������       �        
             2@e      f                    �?��S�ۿ?	             .@������������������������       �؇���X�?             @������������������������       �                      @������������������������       �        	             3@i      n                    �?�R��H�?�           Ј@j      m                   �?�Q���?           �{@k      l                   �?�v�Q�?�            0w@������������������������       ��T��5m�?�             i@������������������������       �N�	g�!�?i            @e@������������������������       �">�֕�?(            �Q@o      p                   �?^�W����?�            v@������������������������       �2S��?H�?q            �e@q      r                   �?��9܂�?i            @f@������������������������       �������??            �Y@������������������������       �v�(��O�?*            �R@t      �                   �?ށ�����?"           d�@u      z                   �?���%�0�?m           ��@v      y                    �?`Ӹ����?!            �F@w      x                   �?ףp=
�?             4@������������������������       �r�q��?	             (@������������������������       �                      @������������������������       �                     9@{      ~                   �?Χ�m�c�?L           x�@|      }                    �?Ʀ-�(��?�             q@������������������������       �fȮ�Б�?I            �_@������������������������       �&���7��?^            `b@      �                    �?:\��M7�?�            �o@�      �                   �?��0u���?K             ^@������������������������       ��w�"w��?.             S@������������������������       �v�X��?             F@�      �                   �?p�ݯ��?Z            �`@������������������������       ����b���?(            �L@������������������������       �P����?2             S@�      �                   �?�g4<��?�           �@�      �                    �?T(y2��?M            �]@�      �                   �?@4և���?             E@������������������������       �ףp=
�?             4@�      �                   �?���7�?             6@������������������������       �                     @������������������������       ��}�+r��?             3@�      �                   �?XI�~�?3            @S@�      �                   �?�C��2(�?             F@������������������������       �$�q-�?            �C@������������������������       �z�G�z�?             @������������������������       �Pa�	�?            �@@�      �                   �?ؓ��M{�?h           0�@�      �                   �?r���"��?�            pv@�      �                    �?��ڂe��?�             r@������������������������       �D������?T            @`@������������������������       ���Q��?d             d@�      �                    �?ꮃG��?6            @Q@������������������������       ��xGZ���?            �A@������������������������       ���.k���?             A@�      �                    �?&>hy���?z            �g@������������������������       �d��4�o�?7            �W@������������������������       ��q�Q�?C             X@�      �                   �?D�C=�}�?�           ��@�      �                   �?����y7�?1           ^�@�      �                   �?��Lɿ��?�           X�@������������������������       �                      @�      �                   �?��Q35��?�           P�@�      �                    �?(N:!���?�           ��@�      �                   �?�J��?�           ��@������������������������       �O)�X�?
           �z@������������������������       �dҁ
_�?�            `q@�      �                   �?��<y�_�?0           p~@������������������������       �(�A����?�             t@������������������������       �<���D�?i            �d@�      �                    �?��_l$�?�            �r@������������������������       ���)�c{�?`             c@������������������������       �(;L]n�?Y            �b@�      �                    �?4S)$&�?�           d�@�      �                   �?p�b孏�?           ��@������������������������       �                     �?�      �                   �?�/���?           ��@�      �                   �?������?N           ��@������������������������       ���Q�`9�?�             w@������������������������       � E�+0+�?c            �c@������������������������       ���S�U�?�            Pr@�      �                   �?�pX�^ѻ?�           ��@�      �                   �?�w��?�           X�@�      �                   �?����y�?           �|@������������������������       �                     @������������������������       �������?           @|@�      �                   �?h�WH��?i            @d@������������������������       �                     @������������������������       �0��_��?h            �c@�      �                   �?�I�R�?           p{@������������������������       �                     @������������������������       ��2c�$��?           0{@�      �                    �?�+�!|�?m           7�@�      �                   �?����	�?�           �@�      �                   �?8ِ��?r           �@�      �                   �?�v�F�?�           ؅@������������������������       �P��k�?+           �|@������������������������       ��J�Yy��?�             n@�      �                   �?��-{��?�            �@������������������������       ��8��8N�?            �@������������������������       �$]^z���?�             m@�      �                   �?��tB��?q           �@������������������������       �xn�-:1�?�            �l@������������������������       ��^l�i��?�           �@�      �                   �?8�G��?�	           `�@�      �                   �?(�ߠ��?i           B�@�      �                   �?����Og�?           ؙ@������������������������       �(?~�Z�?            {@������������������������       �p��Gӹ?�           �@�      �                   �?@ �Z�?[           X�@������������������������       ���g�?�            @k@������������������������       �X���b�?�            u@�      �                   �?0u�����?!           <�@������������������������       ���8�$>�?�            0r@������������������������       ��pK퍅�?c           ��@r  tr  bh�h"h#K �r  h%�r  Rr  (KM�KK�r	  hQ�BP      @B�@    ���@    ���@    �%�@     d�@     ��@    �K�@     t�@     @l@      j@    ���@     0�@     �p@     @o@     @e@     �V@     �d@     �V@      @              Y@     �c@     �X@     �c@       @            �S�@     H�@    ���@     @u@     0u@      ,@     pp@      @     @Z@      @     �Y@      @     �Y@      @     @S@      @      9@                      �?      @             �c@              S@      $@     �L@      "@      :@      "@      8@      "@       @              ?@              3@      �?      @      �?      .@             J�@     `t@     ��@      ^@     ��@     �X@     ܐ@      T@     Ѕ@     �P@     Ѐ@      =@      d@      C@     �w@      *@     �q@      @     �W@       @     �L@      2@      G@      @      &@      (@     ��@      6@     �@      $@     $�@      "@     ��@      �?     ,�@              d@      �?     4�@      (@     ��@      "@     p�@      @     ~@       @     @[@      �?     �@     �i@     ��@     @]@      P@             �@     @]@     ��@     @P@     ��@      J@     L�@     �C@     �p@      *@     X�@     @V@      F@      @      6@      @      6@             ��@     �U@     ��@     �@@     ��@     �J@     8�@     �D@     �i@      (@      h@     ��@      9@      z@      2@     Pu@              *@      2@     �t@      ,@     �f@      ,@     �a@             �D@      @     `b@       @     @Z@       @      E@      @     �R@      @      @@      �?     �E@     �d@     �u@      W@      j@     �J@     �Z@     �C@     �Y@      ;@      S@      (@      :@     �R@     �a@     �P@      ]@      D@     �Q@      :@     �F@      "@      9@     b�@     ��@     ��@     0@     �o@      w@     @a@     �[@      _@     �P@      "@      2@       @      2@      �?             �\@     �H@     �Q@      F@     �H@      F@      6@              F@      @     �D@      @      @              ,@     �E@      @      E@              $@      @      @@      @      �?     �\@     @p@      @      Y@      @     �R@              9@     �[@      d@      X@      [@     �R@     �V@      P@     �V@      &@              5@      1@      2@      1@      @              .@      J@      @      J@       @             ��@      `@      $@             ��@      `@     T�@      I@     �s@      @     �f@      @     �`@             ؆@      G@      �@     �D@     0v@      7@     �k@      2@     `c@      @     ��@     �S@     ��@      M@     �q@       @     �g@      @     @W@      @     ��@      I@     Px@      C@      f@      (@     �k@      5@     �E@      @     @f@      2@      m@     ��@     �^@     І@      @     0�@             �S@      @     p}@       @     �h@      �?      q@     �]@     �f@     �E@      L@      S@      _@     �[@     ��@              8@     �[@     ��@      @     Px@       @     �X@      �?     �A@      �?     �O@      @     0r@      @      \@      �?     `f@      Z@      g@     �C@     @T@      3@      D@      4@     �D@     @P@      Z@      6@     �F@     �E@     �M@     *�@     �@     ��@     M�@     4�@     `�@     <�@     �@     �@      `@     ��@     @P@     �c@     �O@      X@      E@      N@      5@     ��@       @      u@      �?     pr@      �?     �~@     �O@     �Q@      N@      �?      �?     �Q@     �M@      E@     �I@      <@       @     �z@      @     �q@      @     `a@             �x@     �@     �O@     ȅ@      H@     H�@      <@     `i@      4@     �{@      .@      H@      @      6@       @      :@     �t@      $@     �d@      @      \@      @      K@      �?      e@      @     �_@      @      E@             �o@     P}@     @_@     �`@     @T@      9@      ,@      7@     �P@       @      F@     @[@      @     @[@     �B@              `@     �t@      K@      >@      @      >@      H@             �R@     s@      $@     �r@     @P@      @      3@     j�@      (@     ��@      �?     ��@             ��@      �?     @e@      �?      M@              \@      &@     |�@      "@     Ē@      @     �c@      @     P�@       @     �e@             �E@       @     ``@      @     `�@       @     �`@              S@       @     �L@      @     L�@             @|@      @     <�@     �@     ��@     �@     X�@     �@     @p@     Ȓ@     �]@     P�@     �Q@      (@       @      @       @       @             ��@     @Q@     0{@      E@     �p@      ;@     �~@     �G@      x@      C@      @      �?     �w@     �B@     �Y@      "@      @              X@      "@     ��@     �a@      3@      *@      "@       @      @       @      @              $@      &@      @      $@      @      �?     ��@      `@     H�@      J@     @t@      7@     �l@      =@     Py@     @S@     �o@      O@     �b@      .@     �p@     8�@     @V@     �n@     �O@      c@     �B@      R@      :@     @T@      :@      W@      4@     �J@      @     �C@     `f@      w@      b@     �r@      D@     @_@      Z@     `e@     �A@     �R@      *@     �@@      6@     �D@     ؇@     0u@     �q@     �W@     @d@     �G@      a@      0@       @             �`@      0@      :@      ?@      ^@     �G@     �Z@      @      @              Z@      @      *@     �D@     ~@     �n@     �k@     �U@     �e@      0@     �G@     �Q@     0p@     �c@     `i@      @@      @       @     �h@      >@      L@     �_@     .�@     ��@     t�@     ��@     ��@     x�@     ��@     �t@     �y@     `j@       @      4@              *@       @      @      �?      @      �?      @     �y@     �g@     �v@     �f@      j@      Y@      c@     @T@      I@      $@     `s@      ^@      �?             Ps@      ^@     �b@      F@      @      @     @b@      C@     �c@      S@              (@     �c@      P@     �]@      H@     �C@      0@     �~@     @v@      �?     �I@      �?      @@              2@      �?      ,@      �?      @               @              3@     �~@     s@     @q@     �d@     �l@     �a@      `@      R@     �X@     �Q@      H@      6@     �j@     �a@     @\@      O@      Y@     �S@     �L@      G@     �E@      @@      �@     ȁ@      v@     @k@       @     �E@       @      2@       @      $@               @              9@      v@     �e@     �f@      W@     @T@      G@     @Y@      G@     @e@     �T@     �U@      A@     �K@      5@      ?@      *@      U@     �H@      A@      7@      I@      :@     �s@     �u@       @     �[@      @     �C@       @      2@      �?      5@              @      �?      2@      @      R@      @      D@      @      B@      �?      @      �?      @@     `s@      n@     �h@     @d@     @d@      `@      Q@      O@     �W@     �P@     �A@      A@      3@      0@      0@      2@     @\@     �S@      M@     �B@     �K@     �D@     Ѕ@     V�@     @t@     ֧@     @d@     Д@               @     @d@     Ȕ@      a@     x�@     @Q@     Ѓ@     �B@     @x@      @@     �n@     �P@     @z@     �G@     0q@      4@      b@      :@     @q@      5@     ``@      @      b@     @d@     ܚ@     @Y@     ��@              �?     @Y@     ��@     �L@     �}@     �D@     �t@      0@     �a@      F@      o@     �N@     (�@      D@     �@      9@      {@              @      9@     �z@      .@     `b@              @      .@      b@      5@      z@              @      5@     �y@     `w@     ��@     �f@     ��@     �`@     ��@     �G@     `�@      7@     0{@      8@      k@     �U@     ��@     �O@     �@      7@      j@      I@     ��@      *@     @k@     �B@     ��@     �g@     �@      \@     b�@     �T@     ��@      2@      z@     @P@     �@      =@     p�@      .@     `i@      ,@     0t@     �S@      �@      (@     pq@     �P@     ��@r
  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h7Kh8Kh9h"h#K �r  h%�r  Rr  (KK�r  hQ�C              �?r  tr  bhEhUh@C       r  �r  Rr  hYKhZh[Kh"h#K �r  h%�r  Rr  (KK�r  h@�C       r  tr  bK�r  Rr  }r  (hKheM�hfh"h#K �r   h%�r!  Rr"  (KM��r#  hm�Bhk         �                    �?2�Ӛ=��?�e           �@       �                    �?��b���?�5          �@�@       b                    �?�>ٱGx�?�#          �V�@       I                    �?̛��,`�?�          �s�@                           �?p>��5��?G          ���@                           �?����?<           �@                            �?��%�5�?�           P�@                           �?JȬ���?�           ؉@	       
                     �?n9�g���?�           ��@������������������������       ���H��?            |@                           �?����l�?�            `w@������������������������       �dl�'�?�            Pp@                           �?���͡?G            @\@������������������������       �����D��?=            @W@������������������������       �        
             4@������������������������       �                     @                           �?�Y�>3b�?�            �q@                           �?ʐ��7�?�            0q@                           �?$�.Q�,�?�             q@������������������������       �      �?�             n@������������������������       ��������?             A@������������������������       �                     �?                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        �             n@       <                    �?�����ޮ?           �@       -                    �?�[(=�?�           j�@       (                    �?@�k�o��?$           ��@       #                     �?�P��A�?�           ��@                            �?`Ӹ����?           ��@������������������������       �                     �?!       "                    �?��u��ĵ?           ��@������������������������       ���z�Ѻ?\           x�@������������������������       �0;�ø�?�            pr@$       '                    �?B�$U��?�            0u@%       &                    �?�t����?�            �m@������������������������       �                      @������������������������       ��^����?�            �m@������������������������       ���'cy�?E            @Y@)       ,                    �?P��BNֱ?9            �T@*       +                     �?�8��8��?             B@������������������������       �H%u��?             9@������������������������       �                     &@������������������������       �        $            �G@.       5                    �?0g�3c�?�           ׽@/       2                    �?`�j���?�	           ��@0       1                     �?@�f���?           ܟ@������������������������       � b�wKq?�           (�@������������������������       � �#F���?|           h�@3       4                     �?u�6/��?�           ,�@������������������������       � ��h��?�           ܒ@������������������������       ����`�?�           ��@6       9                     �? �*�^�?+	           *�@7       8                    �? �n�EE�?*           ��@������������������������       �        �           <�@������������������������       � U�F.�?U           Ԕ@:       ;                    �?�1��cέ?           D�@������������������������       �        E            �@������������������������       ��_���?�           ��@=       B                    �?�٠n�}�?           ��@>       A                    �?�q�q�?>            �Y@?       @                     �?nM`����?7             W@������������������������       �>���Rp�?"             M@������������������������       �j���� �?             A@������������������������       �                     $@C       F                     �?TK���?�           ��@D       E                    �?��k���?           �z@������������������������       �@�K�҈?w            �d@������������������������       �P#aE�?�            �p@G       H                    �?x�@�E-�?�             t@������������������������       ����1��?A            �Z@������������������������       �Du9iH��?�            �j@J       [                    �?�s_N��?D           ��@K       T                    �?ڵ÷u�?�           ��@L       M                    �?�HK䥲?�            �s@������������������������       �                     .@N       Q                    �?P-�T6��?�            �r@O       P                     �?�߄��i�?�            �l@������������������������       �P���Q�?Z            �a@������������������������       � p�/��?@            @V@R       S                     �? �й���?2            @R@������������������������       �                    �C@������������������������       �г�wY;�?             A@U       X                     �?������?           �y@V       W                    �?��׆�(�?�            �n@������������������������       �8��~P�?S            �^@������������������������       ��4F����?K            �^@Y       Z                    �?�������?n            �d@������������������������       ����3E��?C            @W@������������������������       �P��E��?+             R@\       _                    �?���gb�?f             d@]       ^                     �?�����H�?5            �V@������������������������       �������?            �B@������������������������       ����C��?            �J@`       a                     �?�Y�R_�?1            �Q@������������������������       ��z�G��?             D@������������������������       ��4�����?             ?@c       t                     �?�>`S#�?P           ��@d       o                    �?�#KM�?�           Ж@e       j                    �?܀|��?�           ��@f       i                    �? �Cc}�?             <@g       h                    �?R���Q�?             4@������������������������       ��8��8��?
             (@������������������������       �      �?              @������������������������       �                      @k       n                    �?*`����?�           ؃@l       m                    �?(�\X�?{           �@������������������������       �$��<�?�            `t@������������������������       �����?�            `o@������������������������       ��c�Α�?(             M@p       q                    �?|������?           �@������������������������       ��R����?�            �v@r       s                    �?\�M@��?            {@������������������������       �X�EQ]N�?�             p@������������������������       �&ޏ���?s             f@u       �                    �?�
K5��?�           H�@v       {                    �?<�U����?            {@w       z                    �?@�0�!��?             1@x       y                    �?      �?
             (@������������������������       ��<ݚ�?             "@������������������������       ��q�q�?             @������������������������       �                     @|       }                    �?̠�4��?           �y@������������������������       �D���"�?�            �g@~                           �?~�ו@�?�             l@������������������������       ��Z�K���?m            `e@������������������������       �l��
I��?"             K@�       �                    �?\#r��?{           �@�       �                    �?�*�w�?+            ~@������������������������       �                     �?�       �                    �?Ta'z��?*           ~@������������������������       �ܷ��?��?�            �s@������������������������       �H�ՠ&��?i            @d@�       �                    �?     �?P             `@������������������������       �                     @������������������������       �H�Swe�?O            @_@�       �                    �?��tR��?�           V�@�       �                    �?���SMQ�?           �@������������������������       �                      @�       �                    �?PV�"YP�?           }�@�       �                    �?�Z����?�           ԫ@�       �                    �?�["���?E           Ԡ@�       �                     �?�.7,]�?�            s@�       �                    �?��0u���?p            �f@�       �                    �?4��s?D�?f            �d@������������������������       �N��c��?`            @c@������������������������       ��C��2(�?             &@������������������������       ���S�ۿ?
             .@�       �                    �?��H�}�?G            @_@�       �                    �?�n_Y�K�?A            @]@������������������������       �4uj�w��?=            @\@������������������������       �                     @������������������������       �                      @�       �                     �?�����f�?�           �@�       �                    �?���e��?�           P�@�       �                    �?����պ?           x�@������������������������       ��,/�}�?�            `w@������������������������       �Lq�
���?/           �}@������������������������       ��1=�w��?�            �h@�       �                    �?�����?�           (�@�       �                    �?�!i��?�           ��@������������������������       �`=��?��?�            �p@������������������������       ��~Bo�?�            �v@������������������������       ��E_��?a            �e@�       �                    �?ԳC����?�            �@�       �                    �?L.��:��?C           @@�       �                     �?`׀�:M�?�            �r@������������������������       � ��U��?a            �a@������������������������       ���X8��?g            @c@�       �                     �?�q�q�?{            �i@������������������������       ���Q:��?F            �]@������������������������       �^����?5            �U@�       �                     �?(ڸha!�?@           `�@������������������������       �@�M4��?#            }@������������������������       �0�%�J�?           �{@�       �                    �?��(���?T           &�@�       �                    �?b�u>`�?�           \�@�       �                    �?�ӖF2��?           ��@�       �                     �?���s���?O           ��@�       �                    �?�K�+���?�            Pu@������������������������       ���R[s�?-            �Q@������������������������       �        �            �p@�       �                    �?�:+�X��?t            �g@������������������������       �X�Cc�?             E@������������������������       �@�`%���?\            `b@�       �                    �?C���?�           `�@�       �                     �?z�G�z�?             $@������������������������       �����X�?             @������������������������       �                     @�       �                     �?��p\�?�           �@������������������������       �<�*/�{�?            {@������������������������       ��E�0�/�?�             s@�       �                     �?�kľΣ�?�             k@�       �                    �?�{�@�N�?U            �`@������������������������       �P���Q�?&             N@������������������������       ��1��u�?/            @R@�       �                    �?@4և���?7             U@������������������������       �                     D@������������������������       ���2(&�?             F@�       �                     �?��E�V�?�           ��@�       �                    �?lK��x�?           �y@�       �                    �?�L"p�?f            �d@������������������������       �z�G�z�?             @������������������������       � d�z:�?b             d@������������������������       �xdQ�m��?�            `n@�       �                    �?fRH�w��?�            0r@�       �                    �?���R��?6            @V@������������������������       �                     @������������������������       �v�2t5�?3            �T@������������������������       ���x��?            @i@�       �                    �?�X����?�           \�@�       �                     �?�Ɓ�J�?�            �@�       �                    �?ЋMJ��?           p{@�       �                    �?�<4ޢm�?�            t@�       �                    �?�G�5��?O            @a@������������������������       �>��C��?            �E@������������������������       ��eGk�T�?5            �W@�       �                    �?��GEI_�?w            �f@������������������������       �                     �?������������������������       ����L��?v            �f@�       �                    �?p/3�d��?V            �]@������������������������       ��Fǌ��?6            �S@������������������������       ��e����?             �C@�       �                    �?�#F�\�?�            �t@�       �                    �?���Xr��?�            `j@�       �                    �?�G�z�?             D@������������������������       �����>�?            �B@������������������������       �                     @�       �                    �?�R�+�0�?j            `e@������������������������       �h㱪��?            �K@������������������������       � 	��p�?M             ]@�       �                    �?(��+�?H            �^@������������������������       ���
���?+            �R@������������������������       �p�v>��?            �G@�       �                    �?N�3�t��?�           ��@�       �                    �?�)��V��?f            �d@������������������������       �                     $@�       �                     �?�99lMt�?`            �c@������������������������       �������?0            @U@������������������������       ���U��?0            �Q@�       �                     �?0٘��?S           h�@������������������������       ��7��?�            @m@������������������������       ��IєX�?�            0t@�       p                    �?֚Clb�?0          @��@�       E                   �?�!��?�           �@�       "                   �?�gi��!�?�           �@�       �                    �?��]�Z��?�           �@�       �                    �?D^��#��?            �D@�       �                    �?�ʻ����?             A@�       �                    �?���>4��?             <@������������������������       ����y4F�?             3@������������������������       �                     "@������������������������       �                     @������������������������       �                     @                          �?�nN���?�           l�@                         �?,�x6��?           ��@      	                   �?�����0�?u            `h@                         �?@�k$��?j            �e@                         �?B��仱�?Q            �`@������������������������       ���ꑬ�?D            @[@������������������������       �                     8@                         �?�����?             E@������������������������       �������?            �D@������������������������       �                     �?
                         �?ףp=
�?             4@������������������������       ��t����?	             1@������������������������       �                     @                         �?`����?�           |�@                         �?��l5�̸?0           ��@                         �?��Bb[�?�            0q@������������������������       �0���ަ?r            �e@������������������������       �        B             Y@                         �?@Y.ЂA�?|           X�@������������������������       ���3EaǼ?�             w@������������������������       ��F��O�?�            `k@                         �?B���p�?w             h@������������������������       �tp�P�?D            @[@������������������������       �t�����?3             U@                         �?v���R��?�            �s@                         �?����l�?7            @X@������������������������       � {��e�?            �J@������������������������       �                     F@                         �?�e/
�?�             k@                         �?��.k���?             1@������������������������       ������H�?             "@������������������������       �                      @       !                   �?�`��H �?~            �h@������������������������       �hڛ�ʚ�?`            �b@������������������������       ��+e�X�?             I@#      :                   �?��9���?�           ��@$      /                   �?^+D���?�           ��@%      *                   �?���u��?�            �s@&      '                   �?���ڬ�?�            �p@������������������������       ���n�'��?�            �m@(      )                   �?d��0u��?             >@������������������������       �                      @������������������������       ���2(&�?             6@+      .                   �?�q�q�?             H@,      -                   �?�lg����?            �E@������������������������       ���]�T��?            �D@������������������������       �      �?              @������������������������       �                     @0      5                   �?X@Z@�?�           `�@1      4                   �?�nÈ���?d           Ё@2      3                   �?�������?           0{@������������������������       �        V             a@������������������������       ���ف�"�?�            �r@������������������������       ���7�?\            �`@6      9                   �?�������?�            @n@7      8                   �?`2U0*��?|             i@������������������������       � 7���B�?"             K@������������������������       ����(-�?Z            @b@������������������������       �և���X�?             E@;      @                   �?�����'�?           @}@<      =                   �?�6v��u�?S             a@������������������������       �HQ˄�ľ?C            @[@>      ?                   �?�>4և��?             <@������������������������       �                     �?������������������������       �PN��T'�?             ;@A      D                   �?��B���?�            �t@B      C                   �?�y�b�w�?�             k@������������������������       �                    �B@������������������������       ��,©T�?n            `f@������������������������       ��LQ�1	�?B            �\@F      U                   �?���G��?�           ��@G      L                   �?������?�           X�@H      K                   �?��� �3�?�           8�@I      J                   �?@$��g�?�            �i@������������������������       �                     4@������������������������       ��s0jo�?t            `g@������������������������       �        i           ��@M      P                   �?����h��?�           �@N      O                   �?.�?� ��?�            0q@������������������������       �y�w[��?P            @[@������������������������       ��0���?p            �d@Q      T                   �?T�y���?           ȓ@R      S                   �?�)���Y�?�            �x@������������������������       �                     @������������������������       ��ʈD��?�            0x@������������������������       �ȴ�S뭽?           P�@V      _                   �?XM�N��?            ܢ@W      \                   �?�
��?�           ��@X      Y                   �?p�|�i�?c             c@������������������������       �                     "@Z      [                   �?��LsƔ�?]            �a@������������������������       �                    �E@������������������������       � "��u�??             Y@]      ^                   �?@Vq����?d           0�@������������������������       �        :            �V@������������������������       �`�VX$��?*           �|@`      g                   �?�i�e���?9           ��@a      d                   �?�T_�/��?6           �~@b      c                   �?f1r��g�?�            �j@������������������������       �6�iL�?)            �M@������������������������       �
����?c             c@e      f                   �?�Ug$�Z�?�            Pq@������������������������       ��5��
J�?             G@������������������������       � :��?�            �l@h      k                   �?�G�����?           �@i      j                   �?\X��t�?y            �i@������������������������       �և���X�?&             L@������������������������       ��9��L~�?S            �b@l      o                   �?�.�tT7�?�           ��@m      n                   �?\2R}�?�            r@������������������������       �                     @������������������������       �d�;�s��?�            �q@������������������������       �0w��iv�?�           ��@q      �                   �?r�ܻK�?�           e�@r      �                   �?v�kOSm�?�           y�@s      �                   �?���!���?�           L�@t      �                   �?��z��?           ��@u      |                   �?�O����?�            �q@v      y                   �?���4Z��?�            `p@w      x                   �?P̏����?�            �l@������������������������       ��(\����?4             T@������������������������       ��r*e���?Z            �b@z      {                   �?ҳ�wY;�?             A@������������������������       �                     �?������������������������       ����|���?            �@@}      ~                   �?      �?             6@������������������������       �                     $@      �                   �?�8��8��?             (@������������������������       �؇���X�?             @������������������������       �                     @�      �                   �?�v;�Z�?j           ��@�      �                   �?@B���d�?�           ��@�      �                   �?��<D�m�?Z           ؀@�      �                   �?���N��?h            `c@������������������������       �                     �?������������������������       ��e���@�?g            @c@�      �                   �?8��8���?�             x@������������������������       �                      @������������������������       ��Ht��?�            �w@�      �                   �?0��P�?�            �n@������������������������       �                     �?�      �                   �?��<D�m�?�            �n@������������������������       ��(\����?0             T@������������������������       ���1���?h            �d@�      �                   �?��1[��?w             h@������������������������       ���w/���?Q            ``@������������������������       �V��z4�?&             O@�      �                   �?/]�N��?�           ��@�      �                   �?�	��L��?�           ��@�      �                   �?�(�S	��?`           �@������������������������       ����EƳ?C           @�      �                   �?�Ra����?             F@������������������������       �և���X�?             @������������������������       �@-�_ .�?            �B@�      �                   �?������?�           X�@�      �                   �?�q�w��?,           �}@������������������������       �      �?M             `@������������������������       ���%�r�?�            �u@������������������������       �x���H��?p            �e@�      �                   �?�M���?�             q@�      �                   �?䯦s#�?"            �J@������������������������       �>���Rp�?             =@�      �                   �?r�q��?             8@������������������������       �X�Cc�?             ,@������������������������       ����Q��?             $@�      �                   �?0�й���?�            `k@�      �                   �?`���i��?{             f@������������������������       ������H�?            �F@������������������������       ��	a�$a�?\            ``@������������������������       ��^�����?            �E@�      �                   �?�\Ps��?�
           Ӱ@�      �                   �?���N-�?�           И@�      �                   �? ��&{��?�            �x@������������������������       �        +            �Q@�      �                   �? ��J[�?�            Pt@������������������������       � �IX�-�?�             q@������������������������       ����J��?#            �I@�      �                   �?@�@�{�?�           ��@������������������������       � /��GD?�           P�@������������������������       ��'F�3�?^            �b@�      �                   �?� oA��?�           >�@�      �                   �?���t�?
           x�@�      �                   �?�=��=��?�           0�@������������������������       �                     @�      �                   �?��	��?           �@������������������������       ���7_�?|            �i@������������������������       ��g�y��?           0y@�      �                   �?����?�             m@������������������������       �Z��Yo��?%             O@������������������������       ������?d            `e@�      �                   �?ܾ�z�<�?�           @�@�      �                   �?�_���P�?�             r@������������������������       ��ʹ��Q�?�            �l@������������������������       ��G�z��?$             N@�      �                   �?�y#�Q�?�           ��@������������������������       ��L#���?            ؒ@������������������������       ��	�(�Z�?�            �w@�      �                   �?�\aI5�?           Q�@�      �                   �?�$Ł_�?�           �@�      �                   �?D��?           �{@�      �                   �?؇���X�?F            @Z@�      �                   �?�ʈD��?9            �U@������������������������       �                     4@������������������������       �<���D�?,            �P@�      �                   �?p�ݯ��?             3@������������������������       �                     @������������������������       �        	             (@�      �                   �?PoCFnj�?�            �t@������������������������       ���w�1�?�            r@�      �                   �?*
;&���?             G@������������������������       ��z�G��?             $@������������������������       �                     B@�      �                   �?�6�S2�?�           `�@�      �                   �?hV�a��?d           x�@�      �                   �?�f�¦ζ?G            �Z@������������������������       �0��_��?"            �J@������������������������       �        %             K@�      �                   �?��m�=�?           @|@������������������������       �(���h�?|            �i@������������������������       ��TG!u�?�            �n@�      �                   �?V]��pZ�?b            �c@������������������������       �ƆQ����?(            �N@������������������������       ��q�q��?:             X@�      �                   �?������?*           ��@�      �                   �?��J ��?�           ��@������������������������       �                     @@�      �                   �?��-�=��?�           ��@�      �                   �?b���f�?�             q@������������������������       ������?w             g@������������������������       ���S���?9            �V@������������������������       �� Λ��?           �z@�      �                   �?���ݨ��?O           ޣ@������������������������       � r:�M$p?v           ��@�      �                   �?������?�           �@������������������������       �r�z-��?�            �j@������������������������       ��ę�Z�?T           ��@r$  tr%  bh�h"h#K �r&  h%�r'  Rr(  (KM�KK�r)  hQ�B�      �{�@    ���@    ���@     "�@     L�@     *�@    ���@     ؖ@     6�@     �@     ��@     0}@     �@     0}@     @�@     0s@     (�@     0s@     �m@     `j@     `q@      X@     �d@     �W@     �[@       @     �V@       @      4@              @             @^@      d@      ]@     �c@     �\@     �c@     �V@     �b@      9@      "@      �?              @      �?      @                      �?      n@             }�@      s@    ���@      n@     В@     @R@     ��@     �Q@     ��@      C@      �?             ��@      C@     ��@      ?@      r@      @     0s@      @@     @j@      <@       @              j@      <@     @X@      @      T@      @     �@@      @      6@      @      &@             �G@             /�@      e@     ĭ@      X@     ��@      "@     �@      @     8�@      @     Л@     �U@     �@     �N@     Ѓ@      :@     ��@      R@     B�@     �A@     <�@             H�@     �A@     ��@     �B@      �@             `�@     �B@     ��@     �O@      Q@      A@      M@      A@      F@      ,@      ,@      4@      $@             ��@      =@     z@      *@     `d@      �?     �o@      (@      s@      0@     �Z@      �?      i@      .@     �h@     ��@     �d@     ��@      (@     s@              .@      (@      r@      &@     @k@      @     �`@      @     @U@      �?      R@             �C@      �?     �@@      c@     p@     �U@     �c@     �G@     �R@     �C@      U@     �P@     �X@      C@     �K@      =@     �E@      @@      `@      $@      T@      @     �@@      @     �G@      6@     �H@      (@      <@      $@      5@     8�@     |�@     0�@     p�@     �z@      m@      @      9@      @      1@      �?      &@       @      @               @     �z@     �i@      x@     �g@     �k@     �Z@     �d@     @U@      E@      0@     �U@     0�@      B@     pt@     �I@     �w@      >@     �l@      5@     `c@     v@     ��@     Pr@     `a@      @      ,@      @      "@       @      @      �?       @              @      r@     @_@     `a@     �I@     �b@     �R@     @\@      M@      C@      0@      N@     0�@      K@     �z@              �?      K@     �z@     �@@     �q@      5@     �a@      @     �^@              @      @     �]@     ��@     �@     ȩ@     6�@               @     ȩ@     2�@     ̝@     ܙ@     �@     �v@     �e@     ``@      `@     �I@      `@     �B@     �]@      B@      $@      �?      �?      ,@     �F@      T@     �F@      R@     �D@      R@      @                       @     8�@     `m@     ��@     �]@      �@     �G@     w@      @     �z@      E@     �_@     �Q@     ��@     @]@     X�@     �F@     Pp@       @     `t@     �B@     @Y@      R@     �]@     $�@      R@     �z@      @     @r@      �?     �a@      @     �b@      Q@      a@      F@     �R@      8@      O@     �G@     �@      7@     �{@      8@      z@     ĕ@     �@     �@     `q@     ��@     �V@      @      A@     0t@      2@      J@      2@     �p@             �e@      0@      ;@      .@     @b@      �?     ��@      L@       @       @      @       @      @             `�@      K@      y@      @@     �q@      6@      =@     �g@      7@     �[@      @     �L@      4@     �J@      @     �S@              D@      @      C@      f@     `�@     @[@     �r@     �W@      R@      �?      @     @W@      Q@      .@     �l@     �P@      l@      H@     �D@              @      H@      A@      3@     �f@     (�@     ��@      ~@      r@     @r@     `b@     0q@      G@      Z@      A@      $@     �@@     �W@      �?     `e@      (@      �?             @e@      (@      1@     @Y@      �?     �S@      0@      7@     �g@     �a@     �e@     �B@      *@      ;@      $@      ;@      @              d@      $@     �J@       @      [@       @      0@     �Z@       @     @R@      ,@     �@@     ``@     ��@      Y@     �P@              $@      Y@      L@     �J@      @@     �G@      8@      ?@     p�@      (@     �k@      3@      s@     �@     ��@     J�@     v�@     L�@     ؊@     ��@     �q@      3@      6@      3@      .@      *@      .@      @      .@      "@              @                      @     X�@     Pp@     ��@      h@     @\@     �T@     �[@      P@     @R@      N@     �H@      N@      8@              C@      @     �B@      @      �?               @      2@       @      .@              @     ��@     �[@     ��@      F@     �p@      @     `e@      @      Y@             �@      D@     �u@      6@      i@      2@     �_@     �P@     @R@      B@     �J@      ?@     �n@      Q@     �K@      E@      &@      E@      F@             �g@      :@       @      "@       @      �?               @     �f@      1@      b@      @      C@      (@     �@      �@     h�@     �w@      J@     �p@      B@      m@      9@     �j@      &@      3@       @              @      3@      0@      @@      0@      ;@      .@      :@      �?      �?              @     ȅ@     �\@     ~@     @V@      y@     �@@      a@             �p@     �@@     �S@      L@      k@      :@      h@       @      J@       @     �a@      @      8@      2@      q@     �h@      (@     @_@      @     �Y@      @      7@      �?              @      7@     @p@     �Q@      g@      ?@     �B@             �b@      ?@     �R@      D@     �w@     �@      f@     ��@      @     �@      @     `i@              4@      @     �f@             ��@     �e@     `�@     �T@      h@     �B@      R@      G@      ^@     �V@     `�@      B@     @v@              @      B@     �u@      K@     ��@     �i@     @�@      $@     ��@      @     @b@              "@      @      a@             �E@      @     �W@      @     �@             �V@      @     p|@     �h@     ��@     �I@     `{@      @@     �f@      0@     �E@      0@      a@      3@      p@      &@     �A@       @     �k@      b@     ؐ@     �V@     @]@      8@      @@     �P@     @U@     �K@     �@      4@     �p@              @      4@     �p@     �A@     ��@     Ц@     ��@     �@     x�@     ��@     ��@     ��@     �s@     �S@     �i@      Q@     @h@      L@     �e@       @     �S@      K@     �W@      (@      6@              �?      (@      5@      &@      &@      $@              �?      &@      �?      @              @     (�@     @[@     �@      H@     �@     �@@      c@       @      �?              c@       @     v@      ?@       @             �u@      ?@     �l@      .@      �?             �l@      .@     �S@       @      c@      *@     �`@     �N@     @V@      E@     �E@      3@     ؇@     �@     8�@     �@      9@      �@      4@     �}@      @     �C@      @      @       @     �A@     p�@     @_@     Pz@     �L@      _@      @     �r@     �J@     @Z@      Q@     �j@      N@      4@     �@@      @      6@      *@      &@      "@      @      @      @      h@      ;@     @d@      ,@      D@      @     �^@      "@      >@      *@      u@     �@      &@     ��@      @     px@             �Q@      @     t@      @     �p@      �?      I@      @     ��@      @     @�@      @     @b@     pt@     ��@     @a@     (�@     �Y@      �@              @     �Y@     �@     @V@     �]@      *@     `x@      B@     �h@      7@     �C@      *@     �c@     �g@     L�@     �Y@     `g@      S@     @c@      ;@     �@@     �U@     `�@      R@     ��@      ,@     �v@     8�@     ԫ@     ��@     @     �B@     0y@      .@     �V@       @     �S@              4@       @      M@      @      (@      @                      (@      6@     �s@      .@      q@      @     �C@      @      @              B@     p�@     �W@     (�@      E@     �Y@      @      H@      @      K@             �y@     �B@      h@      *@     �k@      8@     @Z@      J@     �G@      ,@      M@      C@     �j@     �@      R@     ��@              @@      R@     ��@      I@      l@       @     �f@      H@      E@      6@     `y@     �a@     Ƣ@       @     ��@     @a@     ��@      R@     �a@     �P@     ��@r*  tr+  bubhhubh)�r,  }r-  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h7Kh8Kh9h"h#K �r.  h%�r/  Rr0  (KK�r1  hQ�C              �?r2  tr3  bhEhUh@C       r4  �r5  Rr6  hYKhZh[Kh"h#K �r7  h%�r8  Rr9  (KK�r:  h@�C       r;  tr<  bK�r=  Rr>  }r?  (hKheM�hfh"h#K �r@  h%�rA  RrB  (KM��rC  hm�B�d         6                   �?�%�Z���?�e           �@       �                    �?��pp+(�?M:          �-�@                           �?<�O_��?�(           �@                            �?ք:}��?           $�@                            �?�/����?K            �@������������������������       ��j����?           P{@                           �?"� !��?D           �~@                           �?R?4�W�?�            v@	       
                    �?�=~.Y�?�            �u@������������������������       ��1���?�            @n@                           �? '��h�?F            @[@                           �?�f�¦ζ?E            �Z@������������������������       � rpa�?;            @W@������������������������       �        
             ,@������������������������       �                      @������������������������       �                      @������������������������       �        [            �a@                           �?����o��?�            Pr@������������������������       �Ɯ�@Bu�?�            �j@                           �?8�Z$���?3            �S@                           �?�	j*D�?            �C@                           �?p9W��S�?             C@������������������������       �¦	^_�?             ?@������������������������       �����X�?             @������������������������       �                     �?������������������������       �                    �C@       v                    �?>�\�?�%          ���@       ]                    �?������?�           ��@       <                    �?03[�;��?�           �@                           �?���+N�?           ��@������������������������       �                     @        /                    �?�Z���?          ���@!       (                    �?@���z��?3           |�@"       %                     �?XA%�?�           <�@#       $                    �?�}�+r��?           ��@������������������������       � �(�A3�?T           �@������������������������       ��j�j�?�            �p@&       '                    �?ףp=
�?�            �u@������������������������       ��*/�8V�?�            `m@������������������������       ����}<S�?D            �\@)       ,                    �?@�:5�?P	           ڭ@*       +                     �?@�Λۊ?$           ��@������������������������       � ���?           |�@������������������������       ����rݽ�?�           P�@-       .                     �? 8�CS?,           ��@������������������������       �        �           |�@������������������������       � ر��o?:           (�@0       7                    �?���&��?�	           ��@1       4                     �?ؗp�'ʸ?�           ��@2       3                    �?0�C����?�           8�@������������������������       ����7�?             6@������������������������       �������?�           ��@5       6                    �?�b̽s�?�           І@������������������������       �                     2@������������������������       ����M�?�           @�@8       9                    �?�κC��?           b�@������������������������       �                      K@:       ;                     �?��@��?�           �@������������������������       ����w잩?E           ��@������������������������       ���.mZ�?�           x�@=       L                     �?��Hw��?g           L�@>       E                    �?ԣHSp��?u           d�@?       B                    �?V]�t-��?�            �j@@       A                    �?B�~R(��?x            @h@������������������������       ��+��0��?N             `@������������������������       �؇>���?*            @P@C       D                    �?؇���X�?             5@������������������������       ��<ݚ�?             "@������������������������       ��8��8��?             (@F       I                    �?�7,��?�           �@G       H                    �?��P�#��?�           �@������������������������       ���|�r�?�             w@������������������������       �`��4Eѓ?�            0s@J       K                    �?ܢ/��?Q           ��@������������������������       ��p=
�c�?0            ~@������������������������       �<qEH�o�?!           �{@M       N                    �?�ߧ����?�           4�@������������������������       �      �?             @O       V                    �?0�	�t&�?�           �@P       S                    �?�gc� �?�           X�@Q       R                    �?PN��T'�?�            Py@������������������������       ��eP*L��?=            �X@������������������������       ����J��?�             s@T       U                    �?x�}b~|�?�            `u@������������������������       �                     "@������������������������       ��H�@=��?�            �t@W       Z                    �?��j�o�?           �y@X       Y                    �?�q�q�?             �F@������������������������       ��q�q�?            �C@������������������������       ��q�q�?             @[       \                    �?�t��?�            �v@������������������������       ���G^�C�?Z            @`@������������������������       �Dʶ�ˎ�?�            �m@^       m                    �?�=!��M�?N           Ĕ@_       f                     �? �Zz�q�?M           ��@`       c                    �?�뗪K�?�            ps@a       b                    �?Ї���X�?�             l@������������������������       ��t����?             A@������������������������       �@_�M�q�?s            �g@d       e                    �?�6tT�.�?>            �U@������������������������       ��z�G��?             >@������������������������       �0�)AU��?,            �L@g       j                    �?�N8��/�?�            `k@h       i                    �?�9mf��?'            �O@������������������������       ��q�q�?             ;@������������������������       �<ݚ)�?             B@k       l                    �?@f����?^            �c@������������������������       �@�n���??            �Y@������������������������       �                    �J@n       o                    �?�=Z��?           ��@������������������������       �                     *@p       s                     �?�p$orP�?�           ��@q       r                    �?�X�<ݺ?0           @}@������������������������       ������Q�?�            �r@������������������������       ��y��`�?o            �e@t       u                    �?����?�            �s@������������������������       �0�ڂcv�?�            `j@������������������������       � 5x ��?E            �Z@w       �                    �?4N�o;��?�           �@x       �                    �?��-����?�           ��@y       �                    �?4�2%ޑ�?            �A@z       }                     �?����X�?             <@{       |                    �?     ��?             0@������������������������       ������H�?             "@������������������������       �����X�?             @~                           �?�q�q�?             (@������������������������       �և���X�?             @������������������������       ����Q��?             @������������������������       �                     @�       �                    �?R�Ɵ��?�           �@�       �                    �?�p�V��?I           @�@�       �                     �?�^�!<�?S           `�@������������������������       �ʩ�gF%�?�            @u@������������������������       ���.s�?~             k@�       �                     �?�N��?�            �y@������������������������       �    ��?�             p@������������������������       �^Gث3��?c            �c@�       �                     �?�<jV�?L            �^@������������������������       ��GN�z�?)            �P@������������������������       �F�t�K��?#            �L@�       �                     �?/�0r�?           ��@�       �                    �?�Xh�V<�?           �{@������������������������       �                     4@�       �                    �?�H9�^��?           @z@������������������������       �*u�$��?r            �f@�       �                    �?�n\�GZ�?�            �m@������������������������       �ގ$@�h�?g            �c@������������������������       �^�JB=�?8            @T@�       �                    �?\���T��?�            �u@������������������������       �                     :@�       �                    �?�_���?�            @t@�       �                    �?�*|j�#�?�            �o@������������������������       ��fp�I��?h             d@������������������������       ��x�(��?:             W@������������������������       �`��_��?2            �Q@�                          �?��bI���?�           C�@�       �                    �?�ւ�~�?�           ��@�       �                    �?>������?2           X�@�       �                    �?(�� 16�?l            �@�       �                    �?"�����?           �y@�       �                    �?=�Ѝ;�?F            �Y@�       �                     �?�t����?E            �Y@������������������������       �l��
I��?             ;@������������������������       �Х-��ٹ?4            �R@������������������������       �                     �?�       �                    �?BV����?�            ps@�       �                     �?z7Tٲ�?�            �m@������������������������       ����ջ��?F             Z@������������������������       �H�౅z�?T            �`@�       �                     �?؀�:M�?3            �R@������������������������       �������?            �F@������������������������       �П[;U��?             =@�       �                     �?���[�ڥ?Y           0�@�       �                    �? (q~r�?�            0p@�       �                    �?��X8��?i            @c@������������������������       �                     @������������������������       ��'F�3�?e            �b@������������������������       �        @            @Z@�       �                    �?��4+̰�?�            0r@�       �                    �?���%�?u             j@������������������������       �                     �?������������������������       ��R��#�?t            �i@�       �                    �?��`qM|�?;            �T@������������������������       �                      @������������������������       �H�!b	�?:            @T@�       �                    �?�8Ή��?�           ��@�       �                     �?����> �?�           h�@�       �                    �?hu��W�?�             o@������������������������       �,��J�H�?�            @k@������������������������       �r֛w���?             ?@�       �                    �?P���Q�?4           @@������������������������       ����J>�?"            }@������������������������       �@�0�!��?             A@�       �                    �?��H>�6�?�            �w@�       �                     �?�I��쪵?�            �p@������������������������       �p�[&�?Y            �a@������������������������       �     ��?R             `@�       �                     �?@3����?D             [@������������������������       �        #            �K@������������������������       ��&=�w��?!            �J@�       �                    �?*��_��?�           ��@�       �                    �? ,�
-.�?O           �@�       �                    �?&Eȧ��?�           ��@�       �                     �?JJ����?            �G@�       �                    �?��>4և�?             <@������������������������       �                     0@������������������������       ��8��8��?             (@�       �                    �?�d�����?             3@������������������������       �                     @������������������������       ���S�ۿ?
             .@�       �                     �?��
5	�?�           �@�       �                    �?���5��??           �@������������������������       �P�[���?�            �w@������������������������       ��gtq���?N            �`@�       �                    �?�+�cP!�?d           ��@������������������������       �P�19A'�?            z@������������������������       ��M;q��?`            �b@�       �                    �? �-��?�           <�@�       �                     �?�Hy�>d�?�           ��@�       �                    �?���H��?�            `r@������������������������       ������H�?             "@������������������������       �H#���?�            �q@�       �                    �?��`��?�            �v@������������������������       �      �?              @������������������������       �4���?�            pv@�       �                     �?և���X�?�            �w@�       �                    �?�W�,,T�?^             b@������������������������       �����X�?             5@������������������������       ����� �?O             _@�       �                    �?��Ò�[�?�             m@������������������������       � �#�Ѵ�?            �E@������������������������       ��}*��g�?z            �g@�       �                     �?�)p�@�?t            �@�       �                    �?d#����?C           @�@�       �                    �?�\��N��?             3@�       �                    �?ףp=
�?             $@������������������������       �                     @������������������������       �r�q��?             @������������������������       �                     "@�       �                    �?�^����?6           P@�       �                    �?��6L�n�?�            Pt@������������������������       �|�űN�?�            @m@������������������������       �jJA��v�?1            �V@�       �                    �?L���#��?p             f@������������������������       ����C�:�?[            `b@������������������������       �8^s]e�?             =@�       �                    �?    ��?1            �@�       �                    �? �@*��?�            �q@�       �                    �?��<��?~            @i@������������������������       �                     @������������������������       ��ǹ\/�?{            �h@�       �                    �?�	j*D�?(            �S@������������������������       �                     @������������������������       �v���EO�?%            �Q@�                          �?��&y�X�?�             m@                          �?���(`�?e            �e@������������������������       �"pc�
�?             &@������������������������       ��f�?_            `d@                         �?l��[B��?&             M@������������������������       ��q�q�?             @������������������������       ���
ц��?!             J@      !                   �?�������?�           `�@                          �?��Iߪ��?�           ��@                         �?V�a�� �?�            �s@	                         �?��Q��?6             T@
                         �?8�Z$���?            �C@������������������������       �                      @������������������������       ��n`���?             ?@������������������������       �                    �D@                         �?���9yw�?�            �m@                         �?�O2�J�?t             f@������������������������       �؇���X�?             @������������������������       ���Ͻ��?o            @e@                         �?Z��Yo��?)             O@������������������������       �                     "@������������������������       �Ȩ�I��?#            �J@                         �?��1%�?           p{@                         �?ް� ��?B            �Z@                         �?�Zl�i��?3            @T@������������������������       �h�����?             <@������������������������       �^�!~X�?#            �J@                         �?�n_Y�K�?             :@������������������������       �                     $@������������������������       �        
             0@                          �?X�����?�            �t@                         �?@-�_ .�?�            0p@������������������������       ��X�<ݺ?             K@������������������������       ��À���?�            �i@������������������������       ��!�,�E�?+            @R@"      +                    �?��ʃ��?�           ��@#      &                   �?l�R&E�?           �{@$      %                   �?��|.V�?[             b@������������������������       �p���h�?A            @[@������������������������       ��X�<ݺ?             B@'      (                   �?*t�*�N�?�            �r@������������������������       �                     4@)      *                   �?�`K?O��?�            `q@������������������������       ��1j�P�?s            �f@������������������������       ��j&|mH�?=            @X@,      /                   �?�cDh���?�           8�@-      .                   �?LI�#��?�            �u@������������������������       �ܯ/���?�            pq@������������������������       �        (             R@0      3                   �?4և����?�            �x@1      2                   �?��ckݭ�?�            �p@������������������������       �                      @������������������������       �`X�Ɓ5�?�            p@4      5                   �?
XU�)��?S            �_@������������������������       �                     @@������������������������       ����Q��?@            �W@7      �                   �?����N�?=+          @�@8      c                   �?���$���?           B�@9      J                   �?���l��?�           >�@:      A                   �?T���	�?�            �@;      >                    �?�@z�K9�?�            �q@<      =                   �?p����?`             e@������������������������       �                     �?������������������������       �      �?_             e@?      @                   �?���"�?H             ]@������������������������       �                     @������������������������       � '��h�?D            @[@B      E                    �?�L�1�?W           �@C      D                   �?vw۾�+�?T           p�@������������������������       ��c��{-�?W            ``@������������������������       �p#�����?�            �x@F      G                   �?.�	F�9�?           Py@������������������������       �                      @H      I                   �?d�a��M�?           0y@������������������������       ��\�u��?D            �Y@������������������������       ��c��֑�?�            �r@K      \                   �?^!1�I�?�           |�@L      S                    �?H.�!���?             y@M      P                   �?�t%��?�            �k@N      O                   �?�5U��K�?4            �T@������������������������       �                     F@������������������������       �x�����?            �C@Q      R                   �?�I'$;=�?R            �a@������������������������       �~	~���?8            �X@������������������������       ��ՙ/�?             E@T      Y                   �?��]Z�)�?z             f@U      V                   �?Pq�����?:            @U@������������������������       �                     @W      X                   �?������?8            �T@������������������������       ��#-���?            �A@������������������������       �`Ql�R�?            �G@Z      [                   �?n>�X�q�?@             W@������������������������       �*;L]n�?)             N@������������������������       �     ��?             @@]      `                    �? �p�z�?�           x�@^      _                   �?��hwC�?           {@������������������������       ���E�g��?�            �p@������������������������       �Z]k�Β�?h            �d@a      b                   �?d�;�s��?�            �q@������������������������       ���7*��?d            �b@������������������������       ��M8��p�?V             a@d      e                   �?@�O6ٿ�?V           F�@������������������������       �        R            @`@f      w                    �?��!���?           B�@g      r                   �?L��B�?w           �@h      m                   �?���}"c�?P           ��@i      j                   �?(N:!���?�           ��@������������������������       �        x            �g@k      l                   �?h/f���?=           �@������������������������       ����/6��?K            �_@������������������������       ���*>�d�?�            �w@n      q                   �?P� v3t�?�            �n@o      p                   �?�46<�?@             Y@������������������������       ��g�y��?             ?@������������������������       �(���X�?)            @Q@������������������������       ����Hx�?[             b@s      t                   �?\ _;��?'           p}@������������������������       ��Ru߬Α?K            �\@u      v                   �?�����?�            Pv@������������������������       ��2�o�U�?(            �K@������������������������       �I'�2�?�            �r@x      }                   �?���79��?�           h�@y      |                   �?��ٞ?K           X�@z      {                   �?`e	ؚ�?�            pu@������������������������       �`�z�k�?�            �p@������������������������       ��k~X��?,             R@������������������������       �����?�?v            �f@~      �                   �?�"J�?B           <�@      �                   �?.L3�x�?�            �@�      �                   �?~}e}b �?�            �l@������������������������       �2��D�P�?n            `e@������������������������       �Ɣ��Hr�?%            �M@�      �                   �?L�^�?d           ��@������������������������       �x��As�?
           �y@������������������������       �pH����?Z            �`@�      �                   �?�R��(�?K           X�@������������������������       �^%�e��?>            �Z@������������������������       �0�nD-�?           z@�      �                   �?�_E����?          ���@�      �                   �?�n��e��?�	           �@�      �                    �?���̅ӟ?\           Ё@�      �                   �?`#`��k�?�             s@�      �                   �?@�X��?�            `j@������������������������       �@��'��?f             d@������������������������       �p���?             I@������������������������       ��eGk�T�?9            �W@�      �                   �? /8��?�            �p@�      �                   �?�b��fl�?x             g@������������������������       ���<b�ƥ?^            @a@������������������������       �                     G@������������������������       ��(\����?)             T@�      �                   �?�-��>�u?`           ~�@�      �                    �? �&�w]a?�           t�@������������������������       �        �           @�@�      �                   �? d�0�%k?	           Ԓ@������������������������       � �_DT{n?�           Đ@������������������������       �        Z            �`@�      �                    �?�h��4�?�           ��@������������������������       � �[�#�?           �}@������������������������       ��s�k��w?�            �@�      �                   �?�񄔭*�?b           v�@�      �                   �?:9]�w�?X           d�@�      �                   �?�ysT|��?           �{@�      �                   �?�b����?�            u@�      �                    �?dPf�5��?�            �k@������������������������       �6�z���?S            @`@������������������������       ���܂O�?:            �V@�      �                    �?�e"��?N             ]@������������������������       �p�ݯ��?3             S@������������������������       �R���Q�?             D@�      �                    �?l`N���??            �Z@������������������������       �������?!            �O@������������������������       ��^�����?            �E@�      �                   �?xr1�F�?>           ��@�      �                   �? )O��?d            �@�      �                    �?���C:�?            }@������������������������       ����Z�?n            �f@������������������������       �6j\j���?�            �q@�      �                    �?bOvj6��?G            �[@������������������������       �8����?             G@������������������������       �     8�?*             P@�      �                    �?8� WX��?�            �u@������������������������       �bKv���?T            @a@������������������������       �Џxs��?�            �j@�      �                   �?�`�S}�?
           �@�      �                   �?io8�?�	           �@�      �                    �?躘���?�           ƥ@�      �                   �?�Q���#�?	           �@������������������������       � X�}�?           �{@������������������������       ���EOf��?�           ��@�      �                   �?�e�ߧ�?�           ��@������������������������       ���+;Pk�?           �y@������������������������       �x�k6r�?�           ,�@�      �                   �?����p�?�           D�@�      �                    �?���=A��?3           �~@������������������������       �|t���?�            �p@������������������������       �`� x��?�            �l@�      �                    �?0�Ld�?[           �@������������������������       ��w��ݮ?�             l@������������������������       � �b�W�?�            t@�      �                   �?��w�1�?~           R�@�      �                    �?������?P           ��@������������������������       �X�s����?�            �j@������������������������       � ѯ��?�            t@�      �                    �?������?.           (�@������������������������       ��,��v�?�           �@������������������������       ���s�S�?M           D�@rD  trE  bh�h"h#K �rF  h%�rG  RrH  (KM�KK�rI  hQ�B�       ��@     z�@    @6�@     ��@     ��@     ��@     ��@     �|@     ȃ@     �r@     @m@     `i@     �x@      X@     p@      X@     p@     �W@      c@     @V@      Z@      @     �Y@      @      V@      @      ,@               @                       @     �a@             �`@      d@     �P@     �b@     �P@      (@      ;@      (@      ;@      &@      6@      "@      @       @              �?     �C@             <�@     ̔@    ���@     ��@    �v�@     ��@    �(�@     pp@      @             '�@     pp@     �@     @W@     �@     �S@     0�@     �E@     �@      @@     0p@      &@     �s@     �A@     @j@      9@     @Z@      $@     ��@      .@     v�@      ,@     d�@      @     �@       @     ��@      �?     |�@              �@      �?     ^�@     @e@     �@      Y@     h�@      J@      5@      �?     �@     �I@     P�@      H@      2@             ��@      H@     ��@     �Q@      K@             Ԟ@     �Q@     (�@      A@     X�@      B@     8�@     �p@     H�@     �`@     �c@     �L@     �a@      K@     �V@      C@     �H@      0@      2@      @      @       @      &@      �?     З@     �S@     ؄@       @     �v@      @      s@      @     Ȋ@     �Q@     �{@     �@@     �y@     �B@     (�@     ``@      @      @     �@      `@     ��@     �V@     �u@      N@     �F@      K@     �r@      @     �s@      >@      "@             �r@      >@     `w@      C@      >@      .@      :@      *@      @       @     �u@      7@      `@      �?     �j@      6@     (�@     �Y@     @}@      O@     �q@      ;@     `k@      @      >@      @     �g@      �?     @P@      6@      "@      5@      L@      �?      g@     �A@      =@      A@      2@      "@      &@      9@     `c@      �?     �Y@      �?     �J@             ��@     �D@      *@             H�@     �D@     �{@      :@     �q@      &@     �c@      .@     �r@      .@     �h@      (@      Z@      @     �@     ؅@     �@     @v@       @      ;@       @      4@      @      *@      �?       @       @      @      @      @      @      @       @      @              @     Ї@     �t@     Ȅ@     �r@     �x@      d@     �l@     �[@     �d@     �H@     �p@     �a@     �c@     @X@     �[@      G@     @X@      :@     �I@      .@      G@      &@     �{@     pu@     �o@     @g@              4@     �o@     �d@      [@     �R@     @b@      W@      X@     �N@      I@      ?@      h@     �c@              :@      h@     ``@     �c@      X@      X@     @P@     �N@      ?@      B@     �A@     c�@     ��@     >�@     0�@     ��@     H�@      �@     @p@     �d@      o@      *@     �V@      (@     �V@       @      3@      @     �Q@      �?              c@     �c@     �Z@     @`@     �K@     �H@      J@     @T@      G@      <@     �@@      (@      *@      0@     Ѐ@      (@      p@      @     �b@      @      @             @b@      @     @Z@             �q@      "@     `i@      @      �?             @i@      @     �S@      @       @             @S@      @     0z@     (�@      K@     ��@      =@     �k@      5@     �h@       @      7@      9@     �}@      3@     �{@      @      <@     �v@      ,@     0p@      (@     �a@      @     �]@      "@     �Z@       @     �K@             �I@       @     x�@     �@     8�@     �z@     ��@     �e@      6@      9@      1@      &@      0@              �?      &@      @      ,@      @              �?      ,@     0�@     `b@      |@     �O@     �v@      1@     @V@      G@     @~@      U@     �w@      D@     �Z@      F@     ��@     �o@     Ё@     �V@     0p@     �A@       @      �?     `o@      A@     ps@      L@      @      �?      s@     �K@      k@     @d@     �T@      O@      @      .@     @S@     �G@     �`@      Y@       @     �D@     ``@     �M@     p�@     @c@     P|@     �P@      "@      $@      "@      �?      @              @      �?              "@     �{@     �L@     �q@      C@     @k@      0@     @Q@      6@     �c@      3@      a@      $@      4@      "@     �z@     �U@     �m@     �D@      g@      1@      @             �f@      1@      K@      8@              @      K@      1@     @g@      G@     �c@      0@      "@       @     �b@      ,@      <@      >@      @       @      8@      <@     �@     ��@     p�@      i@     �o@     �P@     �G@     �@@      @     �@@               @      @      9@     �D@             �i@     �@@     �d@      $@      @      �?      d@      "@     �C@      7@              "@     �C@      ,@     s@     �`@      2@     @V@       @     @R@      �?      ;@      @      G@      $@      0@      $@                      0@     �q@     �F@     �n@      ,@     �I@      @     @h@      &@      E@      ?@     ��@     `�@     q@     @e@      E@     �Y@       @     @Y@      A@       @     �l@     �P@              4@     �l@     �G@     @d@      3@     @Q@      <@     Px@      v@      V@     pp@      0@     pp@      R@             �r@     �V@     �n@      5@       @             �m@      5@     �L@     �Q@              @@     �L@      C@     ��@     �@     ��@     d�@      x@     t�@     �k@     �@      :@     0p@      5@     �b@              �?      5@     `b@      @     �[@              @      @      Z@     `h@      �@     �[@      z@     �K@      S@     �K@     @u@     @U@      t@               @     @U@     �s@      @@     �Q@     �J@      o@     �d@     Ѝ@      V@     �s@     �I@     �e@       @     �R@              F@       @      ?@     �E@     @X@      ;@     �Q@      0@      :@     �B@     �a@      @     @T@              @      @     �S@      @      @@      �?      G@     �@@     �M@      :@      A@      @      9@     @S@     �@     �L@     �w@      8@     �n@     �@@     ``@      4@     �p@      ,@     �`@      @     ``@     �u@     ��@             @`@     �u@     ��@     �b@     ē@     �\@     �@      T@     `�@             �g@      T@     �z@     �E@      U@     �B@     �u@     �A@      j@      5@     �S@      �?      >@      4@     �H@      ,@     @`@     �A@     @{@      �?     @\@      A@     0t@      1@      C@      1@     �q@     �h@     P�@       @     �@      @     0u@      @     �p@      �?     �Q@      @      f@     �g@     D�@     �`@     �@      X@     �`@     @R@     �X@      7@      B@     �C@     p@      9@     �w@      ,@      ^@     �K@     @}@     �C@     �P@      0@     y@     H�@     S�@      2@     ή@      "@     ��@      @     �r@      @      j@       @     �c@      �?     �H@      �?     �W@      @     0p@      @     �f@      @     �`@              G@       @     �S@      "@     l�@       @     l�@             @�@       @     ̒@       @     ��@             �`@      @     l�@      @     `}@      @     �@     ��@     ?�@     �|@     ��@      c@     0r@      [@     �l@     �Q@     �b@     �J@     @S@      2@     @R@     �B@     �S@      <@      H@      "@      ?@      F@      O@      ?@      @@      *@      >@     s@     h�@     @h@     �w@      c@     �s@      G@     �`@     �Z@     `f@     �D@     @Q@      ,@      @@      ;@     �B@     �[@     �m@      J@     �U@     �M@      c@     �v@     ��@     �l@     �@     �c@     ��@      S@     ��@      3@     �z@     �L@     0�@      T@     d�@      3@     �x@     �N@     8�@     �R@     0�@      G@     |@      =@     �m@      1@     `j@      =@     (�@      @     @k@      6@     �r@     �`@     D�@     �@@     @@      .@     �h@      2@     �r@     �Y@     ��@      9@     P�@     @S@     �@rJ  trK  bubhhubh)�rL  }rM  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h7Kh8Kh9h"h#K �rN  h%�rO  RrP  (KK�rQ  hQ�C              �?rR  trS  bhEhUh@C       rT  �rU  RrV  hYKhZh[Kh"h#K �rW  h%�rX  RrY  (KK�rZ  h@�C       r[  tr\  bK�r]  Rr^  }r_  (hKheM�hfh"h#K �r`  h%�ra  Rrb  (KM��rc  hm�B8i         R                   �?�-�۩��?�e           �@       �                    �?�2�?3E          �@�@       |                    �?<��f�?2          ���@                           �?����B�?�#          �C�@       
                    �?H�z���?h            �@       	                     �?Z`F���?e           ��@                            �?�U�8/��?�           P�@������������������������       ��;�vv��?           `{@������������������������       ����G��?�            @q@������������������������       �z��`p��?�            @n@������������������������       �                     @       A                    �?X���A�?L!          �c�@       2                    �?j!/�H�?�           �@       %                    �?�WG�9��?�           |�@                            �?^��o�?8           ��@                           �?�L���?�           ��@                           �?�U��?e           X�@                           �?�(\����?K             ^@������������������������       �Pa�	�??            �X@������������������������       �                     5@                           �?��Q3��?           ��@������������������������       ��$�'홸?m           �@������������������������       ����Ԋ"�?�            `q@                           �?���BK�?�            �j@������������������������       �����X�?T            �a@������������������������       �x�� ���?/            @R@       "                    �?��9
��?P           �@                           �?|_�,��?�            `w@                           �?��muh�?�            �p@������������������������       ��������?             >@������������������������       �4Q)�i��?�             n@        !                    �?p�eU}�?D            �Y@������������������������       �      �?             @������������������������       � ���v��?@            �X@#       $                    �?4�u���?]            `a@������������������������       ���WV��?E             Z@������������������������       �^������?            �A@&       +                     �?$Q�q�?U            �_@'       *                    �?�?�|�?6            �R@(       )                    �?@4և���?             <@������������������������       ��nkK�?             7@������������������������       �z�G�z�?             @������������������������       �        !             G@,       1                    �?ȵHPS!�?             J@-       0                    �?R���Q�?             D@.       /                    �?����X�?             5@������������������������       �                     �?������������������������       ��z�G��?
             4@������������������������       �        
             3@������������������������       �        
             (@3       :                     �?��
ц��?_            �c@4       9                    �?Hg����?4            �V@5       8                    �?LMc����?.            @T@6       7                    �?���j��?             G@������������������������       �                      @������������������������       �      �?             F@������������������������       �">�֕�?            �A@������������������������       �                     "@;       @                    �?�\����?+            �P@<       ?                    �?V{q֛w�?'             O@=       >                    �?4���C�?            �@@������������������������       �                     �?������������������������       �     ��?             @@������������������������       ��c�Α�?             =@������������������������       �                     @B       a                     �?pl�X�n�?`           ��@C       V                    �?�bV)�X�?u           C�@D       M                    �?0ǹ%�b�?&           ��@E       H                    �?�N�mKs?;           *�@F       G                    �? / �?�           �@������������������������       �        B            �Z@������������������������       ����H��?z           t�@I       J                    �? �3dW?           8�@������������������������       �        "            �M@K       L                    �? ^l� X?]           L�@������������������������       �        �           t�@������������������������       �@t�!�a�?u            �f@N       Q                    �?xD�z�N�?�           �@O       P                    �?�g�%��?�           d�@������������������������       �                     @������������������������       �h֑y��?�           T�@R       U                    �?�oT$?�           l�@S       T                    �?h�����?;            �@������������������������       �                     @������������������������       �0�$<��?8           �@������������������������       ��
#9�?�            0q@W       Z                    �?0�����?O           �@X       Y                    �?h���3}�?           @�@������������������������       �pT[� C�?�            �v@������������������������       �������?#           �{@[       ^                    �?���bXv�?G           ��@\       ]                    �?����X�?�             u@������������������������       �@��,B�?�            q@������������������������       �        ,            �O@_       `                    �?l��\��?v           �@������������������������       �������?           `{@������������������������       ��#-���?\            �a@b       m                    �?B��5��?�	           ��@c       h                    �?@��,B�?H           �@d       g                    �?@or�|ՠ?O           �@e       f                    �?`_U�k-�?�           ��@������������������������       �                     8@������������������������       ������?�           ��@������������������������       ���'����?�            `p@i       j                    �?�4F��?�            �@������������������������       �        {           X�@k       l                    �?�x�V�?~             g@������������������������       �@M^l���?^            �`@������������������������       � ��WV�?              J@n       s                    �?̓��e�?�           �@o       r                    �?�ݩ�v�?~            �@p       q                    �?�`>:��?�           ��@������������������������       �                     @������������������������       �Pd���?�           x�@������������������������       ��� ND��?�            `u@t       y                    �?�G�z�?%            �@u       x                    �?��Ѽ?<           0�@v       w                    �?�܏8o~�?�           h�@������������������������       �                     @������������������������       �ЮN
��?�           0�@������������������������       ����\=y�?�             k@z       {                    �?h�("�?�            �w@������������������������       ��^龆��?�             p@������������������������       �P���Q�?I             ^@}       �                    �?��7�9��?Y           ��@~       �                    �?��w�:��?�           �@       �                    �?��swʭ�?,           `�@�       �                    �?�L�<e�?           x�@�       �                    �?��&�~v�?�           �@�       �                    �?"Xт��?�            �v@�       �                     �?���5��?D            �\@������������������������       ���H�}�?             9@������������������������       ��ƫ�%�?5            @V@�       �                     �?2��8c�?�            �o@������������������������       ��Cc}��?C             \@������������������������       �LRa�v��?]            �a@�       �                     �?xD��t�?�           ��@������������������������       � �P�`��?�            `j@������������������������       �`�q�0ܴ?8           (�@�       �                     �?�9��L~�?g            �b@�       �                    �?L������?7            �S@�       �                    �?r�q��?              E@������������������������       �      �?              @������������������������       �R���Q�?             D@������������������������       �$G$n��?            �B@�       �                    �?*O���?0             R@������������������������       �                     @�       �                    �?h+�v:�?.             Q@������������������������       ���
P��?            �A@������������������������       ����!pc�?            �@@�       �                    �?��Au5a�?           �{@�       �                    �?�t`�4 �?K            �^@�       �                     �?�FVQ&�?            �@@������������������������       �                     @������������������������       ��>����?             ;@�       �                     �?ą%�E�?5            @V@������������������������       ����@��?            �B@������������������������       � pƵHP�?"             J@�       �                     �?�z�G��?�             t@������������������������       �ܾ�z�<�?@             Z@������������������������       � 7���B�?�             k@�       �                    �?�Q�a�~�?�           t�@�       �                     �? ��W�%�?�           ��@�       �                    �?P�4�>�?�            �t@�       �                    �?@�E�x�?z            �h@������������������������       �                     @������������������������       �@��8��?w             h@������������������������       �0�!F��?T            �`@�       �                    �?˒�#�?�            �r@�       �                    �?��Bs�?q            �e@������������������������       �                     @������������������������       �0{�o��?p            @e@������������������������       �4Qi0���?O            �^@�       �                     �?@�?�c�?2           �~@�       �                    �?�J�Է�?�            �n@������������������������       �        \            @b@�       �                    �?@uvI��?<            �X@������������������������       ����J��?!            �I@������������������������       �                    �G@�       �                    �?�g�y��?�             o@�       �                    �?0x�!���?M            �]@�       �                    �?�D�e���?4            @U@������������������������       �                     �?������������������������       ��Ń��̧?3             U@������������������������       ��IєX�?             A@�       �                    �?0Ƭ!sĮ?M             `@������������������������       ��FVQ&�?$            �P@������������������������       �        )            �O@�       �                    �?�AVY��?m           >�@�       �                    �?�����?�           (�@�       �                    �?H5=���?�           @�@������������������������       �                      @�       �                     �?�­v�?�           0�@�       �                    �?�g)k�?�            �x@������������������������       �        	             ,@������������������������       � �qǩ�?�             x@�       �                    �?����p�?           �y@������������������������       �                     @������������������������       ��>����?           Py@�       �                    �?̼Be�z�?�           �@�       �                     �?�J�4�?             9@������������������������       �      �?             (@������������������������       �$�q-�?             *@�       �                     �?TtD9�B�?z           H�@������������������������       ���Fi�1�?�            0p@������������������������       �8��P�?�            `t@�       �                    �?,��S ��?�           T�@�       �                    �?\#r��?!            �N@�       �                    �?�X�<ݺ?             B@������������������������       �                     4@�       �                     �?      �?
             0@������������������������       �      �?              @������������������������       �                      @�       �                     �?�J�4�?             9@�       �                    �?r�q��?             (@������������������������       �z�G�z�?             $@������������������������       �                      @�       �                    �?8�Z$���?             *@������������������������       �      �?             @������������������������       �                     "@�       �                    �?`���i��?�           `�@�       �                     �?0^��2�?�           Ѕ@�       �                    �?�������?�            �v@������������������������       �P���f�?�            �l@������������������������       ��L#���?W            �`@�       �                    �? w���?�            �t@������������������������       ��w��RR�?n            �e@������������������������       �ףp=��?b             d@�       �                     �?e+X�?           ��@�       �                    �?�X��C�?�            �v@������������������������       ��}�+r��?y            �g@������������������������       �XpBt,��?m            �e@�       �                    �? ��<���?           {@������������������������       ��� ND��?{            `e@������������������������       �8Ӈ���?�            `p@�       %                   �? 7�}��?&           �@�                          �?�"�:�I�?/           j�@�       �                    �?&{�7j�?0           h�@�       �                     �?H�!b	�?�            Py@�       �                    �?d��]a��?�            �j@�       �                    �?�w��RR�?i            �e@������������������������       ���*��?T            `a@������������������������       �                    �A@������������������������       ���r._�?            �D@�       �                    �?�eGk�T�?z            �g@�       �                    �?0�)AU��?J            �\@������������������������       �                     "@������������������������       �P�c0"�?E            @Z@������������������������       �        0             S@�       �                     �?:�Q��?5           �}@�       �                    �?��[����?�            Pq@������������������������       ��q�q�?c            �a@�       �                    �?�g+�v�?U             a@������������������������       �r�qG�?@             X@������������������������       �R���Q�?             D@                          �?�y(dD�?}            `h@                         �?(�Z2���?g            `d@������������������������       ��ԇ���?@            �Y@������������������������       ����Q��?'             N@������������������������       �     ��?             @@                          �?P�ihD�?�            �@                         �?�>���?�           H�@                         �?T�6|���?�            �s@������������������������       �                     3@	      
                   �?���ⲣ�?�            Pr@������������������������       �0�z��?�?|            @g@������������������������       �z�H}��?J            �Z@                         �?/8@���?�            s@                         �?H%u��?<             Y@������������������������       �                     F@������������������������       �d}h���?!             L@                         �?��a�Y�?�            �i@������������������������       �                     @                         �?���\��?}            �h@������������������������       �/����?L            �^@������������������������       ��w�"w��?1             S@                         �?�I?YY�?o           ��@                         �?��v����?X           ��@                         �?`��j04�?�            `v@������������������������       �        )             O@������������������������       � c�O�?�            �r@������������������������       �@?�p�?u            @f@      "                   �?p~i��n�?           p|@                         �? i�*$Ŋ?�             s@                         �?@	tbA@�?(            @Q@������������������������       �                     @������������������������       �����e��?'            �P@       !                   �?@���	[�?�            `m@������������������������       �                     8@������������������������       ���^� R�?{            `j@#      $                   �?��)e��?f            �b@������������������������       ��[�IJ�?"            �G@������������������������       �      �?D             Z@&      =                    �?,��ca��?�           3�@'      2                   �?������?�           ̞@(      +                   �?� Luw�?�           �@)      *                   �? ��.lpg?�           Ѕ@������������������������       �@x�5?�?\             b@������������������������       �        a           P�@,      /                   �? �h���?�           ��@-      .                   �? �й���?c            @b@������������������������       ��nkK�?             G@������������������������       �        D             Y@0      1                   �?@p�^5�?c           h�@������������������������       �        /             S@������������������������       ���fh/c�?4           ~@3      8                   �?x���K�?o           Ё@4      7                   �?�Xt��H�?�            `j@5      6                   �?�9ңB��?m            �d@������������������������       ��4�����?@            @W@������������������������       �~X�<��?-             R@������������������������       ��LQ�1	�?             G@9      :                   �?����^��?�            pv@������������������������       �>��C��?r            �e@;      <                   �?vͷu���?q            `g@������������������������       ���S���?            �F@������������������������       ����A��?U            �a@>      G                   �?гY����?            �@?      B                   �?���Ï�?6           `~@@      A                   �?p���ڈ�?�            p@������������������������       � �k/�?d             c@������������������������       �        G             Z@C      D                   �?0�4��?�            �l@������������������������       ��kxipS�?G            @^@E      F                   �?����Z��?D             [@������������������������       �����>4�?!             L@������������������������       �R�}e�.�?#             J@H      O                   �?H��j��?�           4�@I      L                   �?�oY�"T�?�           �@J      K                   �?�P��Э�?<           �@������������������������       � �(�X[o?�           L�@������������������������       ����ƽ�?�             m@M      N                   �?|g�&��?�            `i@������������������������       �        X            �`@������������������������       ���.k���?)             Q@P      Q                   �?�}�+r��?           L�@������������������������       � �(�X[o?�           L�@������������������������       �     8�?{             h@S      �                   �?�^���?�           ���@T                         �?BB!���?�           ��@U      f                   �?�>�u���?�           �@V      e                   �?���Hx�?3             R@W      ^                   �?�y��*�?(             M@X      [                   �?�>4և��?             <@Y      Z                    �?�t����?             1@������������������������       �؇���X�?             @������������������������       �ףp=
�?             $@\      ]                    �?���!pc�?             &@������������������������       �և���X�?             @������������������������       �                     @_      b                   �?��S�ۿ?             >@`      a                    �?@4և���?             ,@������������������������       ��C��2(�?             &@������������������������       �                     @c      d                    �?      �?
             0@������������������������       ������H�?             "@������������������������       �                     @������������������������       �                     ,@g      t                   �?���/6��?{           ț@h      m                   �?m�����?�           l�@i      j                    �?L��f��?]           p�@������������������������       ��G�z��?�             t@k      l                   �?tt���A�?�            �i@������������������������       �                     �?������������������������       ���a�$T�?�            �i@n      q                   �?&�I�f�?M           h�@o      p                    �?�i��M�?�            `y@������������������������       �     .�?�             p@������������������������       ��M;q��?]            �b@r      s                    �?)�p��?R            �]@������������������������       �>���Rp�?(             M@������������������������       ��jTM��?*            �N@u      z                    �?���:�?�           ��@v      y                   �?&RN���?
           @z@w      x                   �?`՟�G��?�            Pu@������������������������       �6�X����?z            �g@������������������������       �z�):���?a            �b@������������������������       ��;u�,a�?/            �S@{      ~                   �?��.b�?�            0s@|      }                   �?��ɍ.�?�            �m@������������������������       �E����?a            `b@������������������������       �n>�X�q�?:             W@������������������������       �j���� �?,             Q@�      �                   �?&�Y����?           0�@�      �                   �?dD�=U�?f           �@�      �                   �?n>�X�q�?           �|@�      �                   �?     ��?             @@�      �                    �?      �?             8@������������������������       �r�q��?             (@������������������������       ��8��8��?
             (@������������������������       �                      @�      �                   �?��J���?�            �z@�      �                    �?330��?�            pq@������������������������       �     ��?K             `@������������������������       ���	c���?Y            �b@�      �                    �?�Ϫ�U�?S            �b@������������������������       ��G�z�?*             T@������������������������       ��û��|�?)            @Q@�      �                    �?D����?Y            �b@�      �                   �?�q�q�?*             R@������������������������       �                     (@������������������������       �z�G�z�?%             N@�      �                   �?"+q��?/            @S@������������������������       �        	             4@������������������������       �F�����?&            �L@�      �                   �?�|�ҵ��?�           X�@�      �                    �?�E����?W            �c@�      �                   �?��a�n`�?              O@������������������������       ��חF�P�?             ?@�      �                   �?�g�y��?             ?@������������������������       �                     "@������������������������       ����7�?             6@�      �                   �?�}�+r��?7            �W@�      �                   �?4և����?!             L@������������������������       ��IєX�?            �I@������������������������       ����Q��?             @������������������������       �                    �C@�      �                   �?��Yז��?^           p�@�      �                    �?��U�I�?�            �p@������������������������       ��P���?J            @\@������������������������       �������?f            �b@�      �                    �?z�RC'��?�            `p@�      �                   �?$��m��?X            @`@������������������������       ��q�q�?              H@������������������������       �H�U?B�?8            �T@�      �                   �?�N2�,��?V            �`@������������������������       ����|���?             F@������������������������       �7�A�0�?9             V@�      �                    �?`�P��˾?�          ���@�      �                   �?TP�m��?�
           (�@�      �                   �?�@t�P�?e           F�@�      �                   �?|n�k�h�?3           ��@�      �                   �?`���pR�?�           8�@������������������������       �                     @�      �                   �?hė+�j�?�           �@������������������������       �p,_�y�?�            @x@������������������������       ���Ջ��?�            �y@�      �                   �?��Ή�ν?5           d�@������������������������       �@-�_ .�?            �{@������������������������       �`�g�ɦ�?           �@�      �                   �?SSx~�?2           �@�      �                   �?�����?           �x@������������������������       �$�q-�?�            @m@������������������������       �XT�z�q�?p            �c@�      �                   �?`�G�Zl�?$           �}@������������������������       ��٠n�}�?�            �n@������������������������       �P���f�?�            �l@�      �                   �?p��*[��?�           �@�      �                   �?     ��?            z@������������������������       �                      @�      �                   �?��g=��?            �y@������������������������       ��חF�P�?[            `c@������������������������       �@-�_ .�?�            0p@�      �                   �?X}�v�?�           (�@������������������������       �\�sl���?�            �j@������������������������       ��y�z���?�           ��@�      �                   �?��@��R�?�           w�@�      �                   �?��`]���?4           x�@������������������������       �                     2@�      �                   �?�ݜۏ��?(           0�@�      �                   �?�t9<��?�           ��@�      �                   �?T�.�"�?�           0�@������������������������       ���� �6�?�            �t@������������������������       �������?           �{@�      �                   �?���b�?�            v@������������������������       ����8��?t            `g@������������������������       �\��1��?d            �d@�      �                   �?��}��?f           (�@������������������������       �T�n��?O             b@������������������������       �0�,���?           P}@�      �                   �? ���*�?�	           2�@�      �                   �?pYnXGG�?           ��@������������������������       �h%Y�b�?           0{@������������������������       �0�>TK�?�           0�@�      �                   �?�}��F̹?�           4�@�      �                   �?��gTj\�?f           ��@������������������������       ���w"�"�?�            �n@������������������������       �Ц�f*�?�            �t@�      �                   �?P�Z��?=           p�@������������������������       ����*�?�            �t@������������������������       �8��O��?|           8�@rd  tre  bh�h"h#K �rf  h%�rg  Rrh  (KM�KK�ri  hQ�B       >�@     ��@    @��@     ��@     ��@     ��@    ���@     ��@     �}@     0~@     �}@     0~@     �x@     �s@     �k@      k@     �e@     �Y@     �S@     �d@      @             �@     ��@     L�@     �r@     ��@      l@     $�@      k@      �@      X@      �@     �C@     @]@      @      X@      @      5@             x�@      B@      �@      =@     �p@      @     �c@     �L@      Y@      D@      L@      1@     �x@      ^@     @t@      I@     `l@      F@      7@      @     �i@     �B@     @X@      @      @      �?     �W@      @     @Q@     �Q@      G@      M@      7@      (@     �]@       @      R@       @      :@       @      6@      �?      @      �?      G@              G@      @      A@      @      .@      @      �?              ,@      @      3@              (@              U@      R@     �J@     �B@      F@     �B@     �@@      *@               @     �@@      &@      &@      8@      "@              ?@     �A@      ;@     �A@      3@      ,@              �?      3@      *@       @      5@      @            ���@     py@     ^�@     �l@     �@      `@     �@      @     �@      @     �Z@             \�@      @     4�@      �?     �M@             H�@      �?     t�@             �f@      �?     ��@     �^@     h�@     �O@      @             X�@     �O@     ��@     �M@     h�@      G@      @             \�@      G@     `p@      *@     X�@      Y@     Ї@      G@     `v@      @     @y@     �C@     ��@      K@     �t@      @     �p@      @     �O@             x�@     �I@     �x@     �C@      `@      (@     .�@     @f@     ��@      3@     h�@      0@     p�@      "@      8@             ��@      "@     �o@      @     �@      @     X�@             �f@      @     �`@      �?      I@       @     Ҡ@     �c@     ��@      S@     0�@      F@      @             �@      F@     `s@      @@     ��@     �T@     ��@      K@     H�@      B@      @             �@      B@     �h@      2@     �u@      =@     `m@      7@     �\@      @     Ư@     Ě@     �@     Ж@     @p@     P�@      m@     ��@     �d@     �@     �^@     �n@      ,@      Y@      "@      0@      @      U@     @[@      b@     �J@     �M@      L@     @U@     �E@     h�@      5@     �g@      6@     �~@     �P@     @U@      D@     �C@     �A@      @      �?      �?      A@      @      @      @@      :@      G@              @      :@      E@      1@      2@      "@      8@      <@     �y@      &@     �[@       @      ?@              @       @      9@      "@      T@       @      =@      �?     �I@      1@     �r@      "@     �W@       @      j@     ��@      @@     Ђ@      7@      t@      "@      h@      @      @             �g@      @      `@      @     �q@      ,@     @e@      @      @             �d@      @      \@      &@     0~@      "@     `n@      �?     @b@             @X@      �?      I@      �?     �G@              n@       @     �\@      @     �T@       @      �?             �T@       @      @@       @     @_@      @      O@      @     �O@             D�@     �o@     (�@      `@     ȇ@     �G@       @             ��@     �G@     �w@      1@      ,@             �v@      1@     �w@      >@      @             pw@      >@     ��@     @T@      5@      @      "@      @      (@      �?     �@     @S@      l@      A@     �q@     �E@     `�@     @_@     �K@      @      A@       @      4@              ,@       @      @       @       @              5@      @      $@       @       @       @       @              &@       @       @       @      "@             ��@     �]@     �@     �L@     u@      ;@     `j@      3@     �_@       @      s@      >@     `d@      &@     �a@      3@      �@      O@     �u@      3@     �f@      $@     �d@      "@     `x@     �E@     `c@      0@     `m@      ;@     (�@     ��@      y@     J�@     `e@     �@      4@     x@      2@     �h@      &@     `d@      &@      `@             �A@      @      A@       @     �g@       @      \@              "@       @     �Y@              S@     �b@     t@     �T@     `h@     �G@     �W@     �A@     @Y@      :@     �Q@      "@      ?@     @Q@     �_@      N@     �Y@      B@     �P@      8@      B@      "@      7@     �l@     ��@     �T@     ��@     �F@     �p@              3@     �F@      o@      @     �f@      E@     @P@      C@     �p@      (@      V@              F@      (@      F@      :@     `f@              @      :@     �e@      @     �]@      5@     �K@     @b@     h�@      R@      }@      @     v@              O@      @     0r@     �P@     �[@     �R@     �w@       @     �r@      �?      Q@              @      �?     @P@      �?     @m@              8@      �?     @j@      R@     �S@      4@      ;@      J@      J@     P{@     ~�@     @h@     ě@      @     ̕@      �?     ȅ@      �?     �a@             P�@      @     Ѕ@       @      b@       @      F@              Y@      @     P�@              S@      @     �}@     �g@     �w@     @P@     @b@     �H@      ]@      >@     �O@      3@     �J@      0@      >@     �^@     �m@      D@     �`@     �T@      Z@      8@      5@     �M@     �T@     `n@     �@     �Q@      z@      @     �o@      @     �b@              Z@     @P@     �d@      D@     @T@      9@     �T@      &@     �F@      ,@      C@     �e@     ڣ@      [@     l�@      S@     ��@       @     D�@     �R@     �c@      @@     `e@             �`@      @@      B@     @P@     H�@       @     D�@     �O@      `@     ֣@     ��@     |�@     ��@     |�@     ؄@      @     @P@      @     �I@      @      7@       @      .@      �?      @      �?      "@      @       @      @      @              @       @      <@      �?      *@      �?      $@              @      �?      .@      �?       @              @              ,@     `�@     Ђ@     ��@     pr@     �x@     �`@     @l@     �W@      e@      C@      �?             �d@      C@     �v@     `d@      q@     �`@     �d@     �V@     �Z@      F@     �V@      =@      F@      ,@      G@      .@     @z@     0s@      m@     �g@     `g@     @c@     �Z@     @U@     @T@     @Q@     �F@      A@     �g@     �]@     �b@     �V@     @V@      M@     �M@     �@@      D@      <@      �@     `�@     `w@     `m@     pr@     �d@      @      =@      @      5@       @      $@      �?      &@               @     @r@      a@     �h@     �T@     @U@     �E@     �[@      D@      X@     �J@      K@      :@      E@      ;@     �S@     �Q@      H@      8@              (@      H@      (@      ?@      G@              4@      ?@      :@     �t@     v@      &@     @b@      @      L@      @      :@      �?      >@              "@      �?      5@      @     �V@      @     �I@      @      H@       @      @             �C@     �s@     �i@     `c@     @[@     �M@      K@      X@     �K@     �d@     �X@     @U@     �F@      @@      0@     �J@      =@     �S@     �J@      <@      0@     �I@     �B@     `�@    ���@     �s@     ܯ@     `l@     ��@     `c@     ��@     �R@     �@              @     �R@     Ȇ@     �A@     v@     �C@     �w@     @T@      �@      8@     @z@     �L@      �@      R@     ؈@     �A@     `v@      2@      k@      1@     �a@     �B@     P{@      2@     @l@      3@     `j@     �U@     ��@     �C@     �w@               @     �C@     pw@      9@     @`@      ,@     �n@      H@     ��@      7@     �g@      9@     ��@      u@     %�@     ``@     l�@              2@     ``@     $�@     �Z@     �@     �R@     ��@     �J@     `q@      5@     `z@      @@     t@      .@     �e@      1@     �b@      9@     `�@      &@     �`@      ,@     p|@     �i@     ��@     �T@     ��@      3@      z@      P@     0�@      _@     <�@      >@      �@      5@     �k@      "@     t@     �W@     ��@      2@     �s@      S@     �@rj  trk  bubhhubh)�rl  }rm  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h7Kh8Kh9h"h#K �rn  h%�ro  Rrp  (KK�rq  hQ�C              �?rr  trs  bhEhUh@C       rt  �ru  Rrv  hYKhZh[Kh"h#K �rw  h%�rx  Rry  (KK�rz  h@�C       r{  tr|  bK�r}  Rr~  }r  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�Bxg         :                   �?������?�e           �@       �                    �?p��k2��?�9          @��@                           �?��q�Y�?"(          @ �@       	                     �?���C���?c           �@                            �?|�{�q�?�           H�@������������������������       ��������?           @z@                           �?8^s]e�?�            Pp@������������������������       �    ���?�             p@������������������������       �                     @
                           �?�����?�             o@������������������������       �ĳ�&���?�            �n@������������������������       �                      @       X                    �?,@~8��?�%          �/�@       1                     �?�5^��?           *�@       &                    �?�LQ�1	�?`           �@       !                    �?��r
'��?#           X�@                           �?����?
           ȓ@                           �?h,H �,�?�           0�@                           �?�2�~w�?�           ��@                           �? �h�7W�?�           ��@������������������������       �h�a��?;            @X@������������������������       ��q�����?a           ؀@������������������������       �      �?	             8@                           �?`Ql�R�?�            �w@                           �?��Y��]�?�            �t@������������������������       �                     *@������������������������       ��u��X�?�            �s@������������������������       �                     H@                            �?��+7��?�            �l@                           �?���!pc�?            �k@������������������������       �������?S             b@������������������������       ���{�?6�?,            �R@������������������������       �                     $@"       #                    �?�8��8��?             B@������������������������       �                     ,@$       %                    �?��2(&�?             6@������������������������       �؇���X�?	             ,@������������������������       �      �?              @'       0                    �?<�;�OK�?=            @Y@(       -                    �?t]����?7            �V@)       ,                    �?���c���?!             J@*       +                    �?��r._�?            �D@������������������������       �                     �?������������������������       �R���Q�?             D@������������������������       �                     &@.       /                    �?�q�q�?            �C@������������������������       ������?             C@������������������������       �                     �?������������������������       �                     $@2       K                    �?:��f	X�?�           Є@3       :                    �?�����?)           }@4       7                    �? �o_��?             9@5       6                    �?z�G�z�?             4@������������������������       ����y4F�?             3@������������������������       �                     �?8       9                    �?���Q��?             @������������������������       �      �?             @������������������������       �                     �?;       F                    �?�7�WR�?           �{@<       C                    �?�>�,M�?�             y@=       @                    �?���@�?�             x@>       ?                    �?0�I��8�?�             o@������������������������       �x��)f��?�            `m@������������������������       �$�q-�?             *@A       B                    �?���.�6�?T            @a@������������������������       �\����?I            @^@������������������������       �                     1@D       E                    �?      �?
             0@������������������������       �؇���X�?             ,@������������������������       �                      @G       J                    �?�\��N��?             C@H       I                    �?����e��?            �@@������������������������       �      �?             :@������������������������       �                     @������������������������       �                     @L       S                    �?7yU�?�             i@M       R                    �?`%za��?a            `c@N       Q                    �?sYi9��?U            `a@O       P                    �?�lhM��?N            �_@������������������������       ��w��d��?:            @W@������������������������       �j���� �?             A@������������������������       �                     (@������������������������       �                     0@T       W                    �?���j��?!             G@U       V                    �?�G�z�?             D@������������������������       �4�2%ޑ�?            �A@������������������������       �                     @������������������������       �                     @Y       �                     �?x��rh��?�            %�@Z       u                    �?�Q��hs�?�           ��@[       h                    �?��@Ԝ~�?�           A�@\       c                    �?�A�tu<�?�	           �@]       ^                    �?@�5|�f�?W           ��@������������������������       �        I            @[@_       b                    �?X�2dgL�?           ��@`       a                    �? ���I�?;           &�@������������������������       ��O"9��?a            �@������������������������       ��@)�<�?�           ,�@������������������������       ����!pc�?�            �t@d       g                    �?܆!+���?�           ��@e       f                    �?0�hz�#�?           (�@������������������������       � qP��B�?�            0x@������������������������       �|�U�7��?(            ~@������������������������       ����e��?o            �h@i       r                    �?(����e�?�           ��@j       m                    �?0�T�5g�?�           |�@k       l                    �? ��R�f?�           ��@������������������������       �        �           x�@������������������������       ����б�?�            �p@n       q                    �?�ƴ�K�?Z           H�@o       p                    �?����Z�?D           �@������������������������       �                     @������������������������       �����)o�?B           ��@������������������������       ��j�+k�?           �|@s       t                    �?�μ���?�            �x@������������������������       �L��G�b�?�            �n@������������������������       �2�6���?]            �b@v                           �?x̓��s�?.           X�@w       |                    �?8��"s�?�           ��@x       y                    �?��S�[�?*            ~@������������������������       �                     @z       {                    �?�d��l��?'           �}@������������������������       �@i�)ԙ�?r            �f@������������������������       ����;QU�?�            @r@}       ~                    �?�{����?�            �o@������������������������       ��Fǌ��?4            �S@������������������������       ���CԐ|�?s            �e@�       �                    �?OX���?]            �a@������������������������       �l��
I��?&             K@������������������������       ��VM�?7            @V@�       �                    �?�X^��B�?�           ��@�       �                    �?x.�[��?           ��@�       �                    �?��@���?�           "�@�       �                    �?WFw:�?6           ��@������������������������       �                     H@�       �                    �?�P�z���?           X�@�       �                    �?��G�ʤ�?4           l�@������������������������       ���&9�J�?�           ��@������������������������       ���(B�@�?�           ��@�       �                    �?�-����?�           D�@������������������������       �        ;           �@������������������������       ����N�.�?�           ��@�       �                    �?(��㓱?�            Ps@������������������������       �        >             Y@������������������������       ��}�+r��?�             j@�       �                    �?
��x�?           �z@������������������������       ��I`Z�?�            �l@�       �                    �?J�8���?�            `i@������������������������       �0N�}S��?c            �c@������������������������       ���+7��?#             G@�       �                    �?X$�`l��?�           x�@�       �                    �?�a:����?,           �@�       �                    �?     7�?�            �@�       �                    �?��z	ÿ?�           H�@������������������������       ��d���?�            Pp@������������������������       � �mѰ��?�            @v@������������������������       �RE��A�?b            �b@�       �                    �?���tT��?C            �@�       �                    �?�|ʉY�?           0z@������������������������       � ��PUp�?Y            �a@������������������������       �	��B�?�            Pq@������������������������       ��E���?B            @X@�       �                    �?,�c�:�?�            @k@�       �                    �?������?e            `d@������������������������       �                     J@������������������������       ��v�ɱ?F            �[@������������������������       �D7�J��?'            �K@�                          �?ʧ"k�E�?�           ��@�       �                    �?08g���?�           *�@�       �                    �?����6W�?�           ��@�       �                    �?&���s�?=           X�@�       �                     �?���C��?A            �Z@�       �                    �?��}*_��?             ;@������������������������       �$��m��?             :@������������������������       �                     �?�       �                    �?pY���D�?.            �S@������������������������       ��g<a�?-            @S@������������������������       �                      @�       �                    �?�W���?�            z@�       �                     �?����i��?�            �s@�       �                    �?��Q�e�?Y             d@�       �                    �?)O���?O             b@������������������������       �p�EG/��?E            �_@������������������������       �        
             2@������������������������       �      �?
             0@�       �                    �?H���I�?c            �c@������������������������       ��q�q�?X            �a@�       �                    �?��.k���?             1@������������������������       �                     @������������������������       �z�G�z�?             $@�       �                    �? %� �?@            �X@�       �                     �?n�C���?:            �V@�       �                    �?*
;&���?             G@������������������������       �r�q��?             E@������������������������       �                     @�       �                    �?F�����?            �F@������������������������       ��s��:��?             C@������������������������       �                     @������������������������       �                      @�       �                    �?����s�?\           ��@�       �                    �?�r��?b           D�@������������������������       �                     1@�       �                     �? ^6�ι?W            �@�       �                    �?Pgi��D�?>           (�@�       �                    �?���J��?�            �o@������������������������       �������?q            �e@������������������������       �        <            �T@�       �                    �?�IєX�?�           0�@������������������������       �8	A�"�?�            y@������������������������       ����X=P�?�            �n@�       �                    �?��Rꉼ?           ؉@�       �                    �?�C͑V�?�            �o@������������������������       �`<�Gf�?q             e@������������������������       � qP��B�?6            �U@�       �                    �?���ÿj�?r           ��@������������������������       �TC��3��?�            `x@������������������������       ���E�"�?u            �f@�       �                     �?��j\���?�             x@�       �                    �?*jF���?o            `d@������������������������       ��^�����?C            �U@������������������������       �:���u��?,            @S@�       �                    �?j@ �'��?�            �k@������������������������       ����p9W�?]             c@������������������������       ��J�T�?.            �Q@�       �                    �?���?#           ��@�       �                    �?���'���?�           �@�       �                     �?H"���?�           ؇@�       �                    �?r�q��?�             n@������������������������       �(N:!���?�            @j@�       �                    �?��S���?             >@������������������������       �                     ,@������������������������       �      �?             0@�       �                    �?�!�d�к?:           X�@������������������������       �%Xhqv�?           �}@�       �                    �?"pc�
�?             F@������������������������       ��eP*L��?             &@������������������������       ��FVQ&�?            �@@�       �                    �?�iZE��?�           0�@�       �                    �?��<��C�?3           ��@�       �                     �?P�H�}��?�            �m@������������������������       ��Ń��̧?M            �_@������������������������       � \sF��?L            @\@�       �                     �?�l���?�           8�@������������������������       �p#x��?�            �r@������������������������       �󝢸]�?�            �u@�       �                     �?�'�^�2�?�            `q@������������������������       ��f7�z�?O             ]@������������������������       ����3L�?k            @d@�                           �?��5bh�?]           (�@�                          �?>ߗ6���?�            �r@�       �                    �?4Q)�i��?�             n@�       �                    �?��It��?2            �S@������������������������       ��z�G��?             >@������������������������       �@�E�x�?            �H@�                           �?h�WH��?]            @d@������������������������       �ףp=
�?             $@������������������������       �@݈g>h�?V             c@                         �?h�����?              L@������������������������       �                     $@������������������������       �(옄��?             G@      
                   �?x��HF�?�            �q@                         �?\�Uo��?             C@������������������������       �d}h���?             <@      	                   �?ףp=
�?             $@������������������������       �z�G�z�?             @������������������������       �                     @                         �?�DS�B�?�            �n@                         �?|_�,��?t            `g@������������������������       ��ʈD��?            �E@������������������������       �8��8���?[             b@������������������������       �TV����?"            �M@      !                   �?*�ߜ�?�           8�@                          �?�q�q�?�           �@                         �?6��h'�?�            �n@                         �?���(\O�?g             d@������������������������       �                      @                         �?�˹�m�?`             c@������������������������       ���E�B��?            �G@������������������������       �T>D5j�?E            @Z@������������������������       �        ,            �U@                         �?(	[\�c�?0           �~@������������������������       �                     =@                         �?��#N�R�?           �|@                         �?\�sե��?H            �\@������������������������       ���IF�E�?%            �P@������������������������       �@9G��?#            �H@                          �?���]�?�            �u@������������������������       �(YB���?�            �p@������������������������       ��Fǌ��?*            �S@"      /                   �?� V�*�?           ��@#      (                   �?�f�?           x�@$      '                    �?r�q��?             2@%      &                   �?      �?             (@������������������������       ����!pc�?             &@������������������������       �                     �?������������������������       �                     @)      ,                   �?�<x�(��?�           �@*      +                    �?���7�?�             v@������������������������       �x�{�;��?f             e@������������������������       �8��"s�?p            �f@-      .                    �?0�E��?(           �{@������������������������       � .2��A�?|            �g@������������������������       �����?�            p@0      5                    �?�!�;��?           �{@1      2                   �?�[�IJ�?u            �g@������������������������       �                    �@@3      4                   �?��`f8�?_            `c@������������������������       �������?$             N@������������������������       �V���#�?;            �W@6      7                   �?Hj�́/�?�            p@������������������������       �        $            �P@8      9                   �?�c)�s�?t            �g@������������������������       ����Q��?3            @U@������������������������       ��k��V��?A            �Z@;      �                   �?�*/���?�+          �;�@<      k                   �?�YՁ�j�?           ��@=      T                    �?�q�!�Y�?�           ��@>      M                   �?P� �&�?�           ��@?      F                   �?x�t�Ap�?           p�@@      C                   �?�zvܰ?�             v@A      B                   �?ps��pй?l             e@������������������������       ��	a�$a�?U            ``@������������������������       �                     C@D      E                   �?��v$���?z            �f@������������������������       �     ��?X             `@������������������������       � �Jj�G�?"            �K@G      J                   �?:ɨ��?           �|@H      I                   �?    �O�?�             p@������������������������       ��?C���?`            �c@������������������������       � %� �?A            �X@K      L                   �?�_�Q��?{            �i@������������������������       �4V��X�?T            `a@������������������������       �P�~D&�?'            �P@N      Q                   �?�rL+��?�            �h@O      P                   �?��v����?-            �P@������������������������       �ܷ��?��?             =@������������������������       ��S����?             C@R      S                   �?&^�)b�?T             `@������������������������       �        4            �S@������������������������       ���.k���?             �I@U      `                   �?�ޡlpg�?'           ��@V      ]                   �?qАݙ�?           �|@W      X                   �? E59|�?~             h@������������������������       �                     &@Y      Z                   �? ��WV�?x            �f@������������������������       �@��8��?A             X@[      \                   �?���1j	�?7            �U@������������������������       ��IєX�?             A@������������������������       �0G���ջ?!             J@^      _                   �? 
�V�?�            �p@������������������������       ��NM�g�?`            �e@������������������������       �        A            �W@a      f                   �?P��e��?           @z@b      e                   �?�~Np���?�            �k@c      d                   �?�M�E$g�?p            �g@������������������������       ��As`�?D            �[@������������������������       �*-ڋ�p�?,            @S@������������������������       �����X�?            �A@g      j                   �?��;���?�            �h@h      i                   �?�I�w�"�?a             c@������������������������       �d,���O�?C            �Y@������������������������       �z�G�z�?             I@������������������������       ��q�q�?             �F@l      w                    �?x:�U��?k           H�@m      r                   �?���l'��?           t�@n      o                   �?      �?           ��@������������������������       ��?�P�a�?�            �v@p      q                   �?x�5?,R�?            {@������������������������       �`RC4%�?�             q@������������������������       �      �?k             d@s      t                   �?Z���t�?x           (�@������������������������       �����^��?8           �}@u      v                   �?|E+�	��?@           `~@������������������������       �����?�            Pp@������������������������       �HP�s��?�             l@x      �                   �?����?�           �@y      ~                   �?�:�1��?�           @�@z      }                   �?  6�W �?,           �}@{      |                   �?p���A�?�             r@������������������������       �                     @������������������������       �ę��N��?�            �q@������������������������       �p�/E�f�?v            �g@      �                   �?4J��4�?�           ��@������������������������       �І�^���?           �|@������������������������       �|�9ǣ�?�            �m@�      �                   �?�I�R�?           p{@������������������������       � �#�Ѵ�?S             `@������������������������       �Hn�.P��?�            `s@�      �                    �?��u#�?�           4�@�      �                   �?\g5�s��?�           ܲ@�      �                   �?t`��q�?.           �@�      �                   �?�3�ڕ?D           ��@�      �                   �?���b��?�            �m@�      �                   �?0���{�?z            �i@������������������������       �                     5@������������������������       �p��ӵ6�?k            �f@������������������������       �                     A@�      �                   �?�]�-/��?�           ��@������������������������       � "�^�?n           ��@������������������������       �        A             X@�      �                   �?hN�����?�           h�@�      �                   �?�Xbv���?�           `�@������������������������       �                     @�      �                   �?2~^�8��?�           H�@�      �                   �?�{%ِ��?;           @������������������������       �>�Q��?H             Z@������������������������       �HX���?�            �x@�      �                   �?6�`��V�?�             o@������������������������       �|�U&k�?*            �R@������������������������       �󝢸]�?k            �e@�      �                   �?�j�-��?           ��@�      �                   �?^��e��?�            �j@������������������������       ��T`�[k�?h            �c@������������������������       �����0�?             K@�      �                   �?���xr�?�           d�@������������������������       �pݲ��l�?�           8�@������������������������       �X	
bi��?�            @n@�      �                   �?y�̆��?�           ��@�      �                   �?��p��P�?B           ؀@������������������������       �                     .@�      �                   �? �	.��?:           `�@�      �                   �?T���ʴ�?|            �h@������������������������       �(;L]n�?M             ^@������������������������       �t�C�#��?/            �S@������������������������       �p���.�?�            Pt@�      �                   �?�QF+�?_            �@������������������������       �                   �{@�      �                   �?���DPF�?F           x�@������������������������       ��_��_�?\            �a@������������������������       �0h�7��?�           �@�      �                   �?Ȓ�g;�?�           ��@�      �                   �?(�Y�$��?�
           ��@�      �                   �?$�А���?           ��@�      �                   �?� ����?           py@������������������������       �        (             O@�      �                   �?�]���?�            �u@������������������������       �0l9i�?�            `r@������������������������       ����J��?&            �I@�      �                   �?�Ha-��?           x�@�      �                   �?JP�ؓ�?�           �@������������������������       ��JY�8��?p             i@�      �                   �?���g�X�?&           �{@������������������������       �                      @������������������������       �h4�)�u�?$           p{@�      �                   �?Hя8X8�?�            �i@������������������������       �θ	j*�?"             J@������������������������       ��s�c���?d            @c@�      �                   �?$�p#�?�           ��@�      �                   �?���/�u�?�           @�@������������������������       ����bȸw?�           $�@������������������������       �`��(�?Z            �`@�      �                   �?LL�lG��?�            �@�      �                   �?$�jkq�?�            �t@������������������������       ��T��5m�?�            �p@������������������������       ��-ῃ�?*            �N@�      �                   �?���s��?�           ��@������������������������       ��^�;��?           |�@������������������������       ��X�<ݺ?�             r@�      �                   �? A��JJ�?7           ��@�      �                   �? YyH9�?           ��@�      �                   �?0�,���?             i@������������������������       �                     <@������������������������       �Ѝܯ0$�?p            �e@������������������������       ����%�<p?�           x�@�      �                   �?4uUD�>�?(           ,�@�      �                   �?��B�5��?D           0�@������������������������       ��q�q�?B             [@�      �                   �?P�cZY�?           �y@������������������������       �                     @������������������������       ��W2ٖ�?�            Py@�      �                   �?`�r�g��?�           @�@������������������������       �:�w�9o�?�            �k@������������������������       ��?�C<�?X           Ĕ@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B�      �o�@    ���@    @��@     X�@    �o�@     ��@     �~@     �{@     �x@     �q@      k@     `i@     �f@     @T@     �e@     @T@      @             �V@     �c@     @V@     �c@       @            �{�@     ��@     t�@     �w@     �@     �f@     (�@     �a@     �@     �Z@     �@     �G@     h�@     �C@     ��@      B@      W@      @     �@      ?@      5@      @      w@       @      t@       @      *@             0s@       @      H@             @e@      N@      d@      N@      Z@     �D@      L@      3@      $@              @     �@@              ,@      @      3@       @      (@      �?      @      M@     �E@      M@     �@@     �F@      @      A@      @              �?      A@      @      &@              *@      :@      (@      :@      �?                      $@     �}@      h@     0x@     �S@      2@      @      0@      @      .@      @      �?               @      @       @       @              �?     w@     �Q@     �u@     �J@     �u@     �C@     @k@      >@     �i@      =@      (@      �?      `@      "@      \@      "@      1@               @      ,@       @      (@               @      4@      2@      4@      *@      *@      *@      @                      @     �U@     �\@     @R@     �T@     @R@     �P@     �N@     �P@     �D@      J@      4@      ,@      (@                      0@      *@     �@@      *@      ;@       @      ;@      @                      @     -�@     ��@     Y�@     ��@     C�@     �@     ��@     `q@     X�@     �c@     @[@             ~�@     �c@     ��@      Q@      �@       @     <�@      N@      n@     �V@     ��@      ^@     ��@     �F@     �w@      "@     �{@      B@     �^@     �R@     Ȫ@      m@     �@     @R@     ��@       @     x�@             �p@       @     ,�@     �Q@     x�@     �B@      @             h�@     �B@     �z@      A@     �m@     �c@     �d@     �T@     �R@     @S@     ��@     @U@     ��@      D@     �|@      7@      @             0|@      7@     `f@      @      q@      4@     `m@      1@     �S@      �?     �c@      0@     �X@     �F@      C@      0@      N@      =@     �@     �y@     ڧ@     `j@     ��@      T@     .�@     @Q@      H@             ΢@     @Q@     Г@     �C@     ��@      @     ��@      @@     ̑@      >@     �@             ��@      >@     �r@      &@      Y@             �h@      &@     �r@     ``@     �d@     �N@     �`@     �Q@     �X@      M@      A@      (@     P�@     @i@     d�@     `e@     ��@     @Z@      �@     �D@     �o@      @     t@     �A@     �U@      P@      |@     �P@     Px@      >@     �a@       @      o@      <@     �N@      B@     `g@      ?@     �c@      @      J@             �Z@      @      <@      ;@     ²@     l�@     �@     |�@     ��@     p�@     �i@     �s@      (@     �W@      $@      1@      "@      1@      �?               @     @S@       @     �R@               @      h@      l@     @_@      h@     @Q@     �V@      Q@      S@      I@      S@      2@              �?      .@      L@     �Y@     �G@     �W@      "@       @      @               @       @     �P@      @@     �P@      8@     �C@      @     �A@      @      @              <@      1@      5@      1@      @                       @     �@     �i@     ԙ@      W@      1@             ��@      W@     Њ@     �E@     @o@      @     �d@      @     �T@              �@      C@     �w@      3@     @l@      3@     P�@     �H@      o@      @     �d@      @      U@       @     ��@      E@     pv@      ?@     `e@      &@     �p@     �\@     �]@     �F@      N@      :@      M@      3@      c@     �Q@     @Z@     �G@      H@      7@     �@     D�@     ,�@     ��@     @Q@     ��@      D@      i@      8@     @g@      0@      ,@      ,@               @      ,@      =@     �~@      5@     �|@       @      B@      @      @       @      ?@     0�@     �h@     (�@     @T@     �l@       @     �^@      @      [@      @     ��@     @R@      q@      ;@     �r@      G@      d@     @]@      Q@      H@     @W@     @Q@      {@     �b@     �l@      Q@     �i@     �B@     �L@      6@      "@      5@      H@      �?     `b@      .@      "@      �?     @a@      ,@      9@      ?@              $@      9@      5@     `i@     @T@      .@      7@      @      6@      "@      �?      @      �?      @             �g@      M@     @d@      9@     �C@      @     �^@      5@      :@     �@@     ܒ@     ��@     �n@     �~@     �Y@     �a@      1@     �a@               @      1@     �`@      @     �D@      &@     �W@     �U@             �a@     �u@              =@     �a@      t@      K@     �N@      @     �M@     �G@       @     @V@     0p@      &@      p@     �S@      �?     �@     �r@     H�@     �Q@      .@      @      "@      @       @      @      �?              @             І@     �P@      u@      0@     `d@      @     �e@      $@     �x@     �I@      e@      3@      l@      @@      k@     �l@      [@      T@             �@@      [@     �G@      F@      0@      P@      ?@      [@     �b@             �P@      [@     �T@     �I@      A@     �L@     �H@     t�@     i�@     0�@     !�@     �t@     l�@      g@     ȉ@      c@     ��@      (@     @u@      "@      d@      "@     �^@              C@      @     �f@       @     �_@      �?      K@     �a@      t@     �S@      f@     �G@     �[@      @@     �P@     �N@      b@     �E@      X@      2@     �H@     �@@     `d@      "@      M@      @      :@      @      @@      8@     @Z@             �S@      8@      ;@     �a@     �@      "@     @|@      @     @g@              &@      @     �e@       @     �W@      @     @T@       @      @@      @     �H@       @     �p@       @     `e@             �W@     �`@     �q@     �T@     �a@     @R@     �\@     �E@      Q@      >@     �G@      $@      9@     �I@     @b@      B@      ]@      :@      S@      $@      D@      .@      >@     �q@     �@     �c@     �@     �X@     ��@      E@     �s@     �L@     pw@     �B@     `m@      4@     �a@     �L@     `�@      2@     �|@     �C@     �{@      5@      n@      2@     �i@     @`@     �@     @[@     ��@      O@     �y@     �D@     �n@              @     �D@     `n@      5@     �d@     �G@     (�@      9@     �z@      6@     �j@      5@      z@      @     �^@      .@     pr@     ��@    �X�@      y@     J�@     �p@     Ԥ@      $@     ��@      @      m@      @     �h@              5@      @     @f@              A@      @     `�@      @     `�@              X@     Pp@     T�@      _@     ��@              @      _@     h�@     �S@     0z@     �@@     �Q@     �F@     �u@      G@     @i@      7@     �I@      7@     �b@      a@     ��@     �K@     �c@      B@     �^@      3@     �A@     �T@     8�@     �O@     @�@      3@     �k@     ``@     ��@      J@     p~@              .@      J@     �}@     �@@     �d@      @      ]@      =@      I@      3@      s@     �S@     �@             �{@     �S@      �@     �K@     �U@      8@     H�@     (�@     g�@     `u@     Ю@      a@     t�@      @     y@              O@      @     0u@      @     r@      �?      I@     ``@     `�@     �X@     ��@     �R@     �_@      8@     z@               @      8@     �y@     �@@     �e@      1@     �A@      0@     @a@     �i@     �@      @     ,�@      @     �@       @     �`@      i@      �@     �]@     `j@      X@     �e@      6@     �C@     �T@     ��@     �P@     t�@      0@      q@     �i@     ��@       @     ��@      @     `h@              <@      @     �d@       @     h�@     �h@     <�@      O@     �|@     �F@     �O@      1@     �x@              @      1@     @x@      a@     �@     @P@     �c@      R@     ��@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�Bxg         J                   �?�J����?�e           �@       �                    �?��E>iJ�?rM          @��@       �                    �?��]�0�?�1          ���@                           �?Ȕ���?�$           %�@                           �?��d:��?s           �@                           �?�=^��?q           ؏@       
                     �?������?n           ��@       	                     �?TB�f�:�?�           ��@������������������������       ��|v���?(           �}@������������������������       ��q�q��?�             r@������������������������       ���8�ͻ�?�             o@������������������������       �                     @������������������������       �                      @       Q                    �?\�8����?S"          �&�@       @                    �?�Oˉۼ�?l           �@       -                    �?0VJr@�?�           $�@                            �?�,f�pY�?           ��@                            �?{�
;�?�           @�@                           �?��arO�?I           ��@                           �?�d���?{            �e@������������������������       ��}�+r��?7             S@������������������������       �        D            �X@                           �?�ɮ�D��?�           |�@������������������������       ���U�(�?a           ��@������������������������       ��u1 e��?m           ��@                           �?��}S߷?Y           ��@                           �?��ϭ�*�?$             M@������������������������       ����N8�?             5@������������������������       �                    �B@                           �?����ɶ?5           Ȍ@������������������������       � ��P0�?�            �o@������������������������       �0v��ꛠ?�           ؄@!       &                     �?`GN6s�?z           �@"       #                    �? �
��>�?�           d�@������������������������       �        (            �N@$       %                    �? >��@�?�           p�@������������������������       �@9G��?�            `r@������������������������       �                   ؒ@'       *                    �?�x��e�?�           ��@(       )                    �?���7�?             6@������������������������       �z�G�z�?             @������������������������       �        
             1@+       ,                    �? ��eҢ�?�           ��@������������������������       ��o�s(��?G            �[@������������������������       �����!sp?D           @.       9                     �?��ș�&�?�	           4�@/       4                    �?�2�{�е?n           R�@0       1                    �?�h[�뱺?�           ��@������������������������       �                     @2       3                    �?����̺?�           ��@������������������������       ��LQ�1	�?             7@������������������������       ���Rqy �?�           @�@5       6                    �?�z�|��?u           ��@������������������������       �                     @@7       8                    �?��¬_��?_           t�@������������������������       �                     @������������������������       ����}�
�?[           \�@:       ;                    �?��\̭ƶ?g           ĕ@������������������������       �                      @<       =                    �?�f�¦ζ?e           ��@������������������������       �                    �B@>       ?                    �?�x�*f�?O           (�@������������������������       ��M8��p�?�           h�@������������������������       �hd�)�b�?�           �@A       J                    �?�Y�R_�?{           �@B       E                    �?�j&|mH�?h           0�@C       D                     �?�+e�X�?             9@������������������������       ��<ݚ�?
             2@������������������������       �����X�?             @F       G                     �?�J����?Y           h�@������������������������       ����W$��?�            �s@H       I                    �?��^@t�?�             n@������������������������       �                      @������������������������       �h�w��?�            �m@K       N                    �?����?           �y@L       M                     �?؇���X�?	             ,@������������������������       �ףp=
�?             $@������������������������       �      �?             @O       P                     �?��D�3��?
           �x@������������������������       ���˙�
�?�            @o@������������������������       ������?h            �b@R       q                    �?4�U>���?�           F�@S       b                     �?p��'���?,           �@T       [                    �?�䳿I��?R           ��@U       X                    �?*��r��?�            �n@V       W                    �?<��u�?�            �l@������������������������       �f�Sa6T�?S            @b@������������������������       �r�q��?2             U@Y       Z                    �?�IєX�?	             1@������������������������       �ףp=
�?             $@������������������������       �                     @\       _                    �? p�۹?�           �@]       ^                    �?����?}           ��@������������������������       ��u��Ek�?�            pu@������������������������       �`��>�ϗ?�            �o@`       a                    �?h�1ڱ��?G           X�@������������������������       ��ꪚ<
�?%           P~@������������������������       ���ӵ�)�?"           `|@c       j                    �?�C��2(�?�           ��@d       g                    �?̚f��p�?]           ��@e       f                    �?��cɻ�?�            �v@������������������������       ��q�Q�??             X@������������������������       �8M��ap�?�            �p@h       i                    �?��A9G�?v            �h@������������������������       �և���X�?            �A@������������������������       �@��'��?a             d@k       n                    �?hz$|b��?}           (�@l       m                    �?���Zdt�?�            @t@������������������������       ��IєX�?             1@������������������������       �0�>TK�?�            0s@o       p                    �?��1���?�            p@������������������������       �                     @������������������������       �����y7�?�            @o@r       y                     �?��D)4�?�           ��@s       v                    �?2G���U�?            z@t       u                    �?��2(&�?             6@������������������������       �ףp=
�?             $@������������������������       �r�q��?             (@w       x                    �?��	t1��?�            �x@������������������������       ��!ݣ�-�?�            �l@������������������������       �����+�?j            `d@z       }                    �?�!���?�            0q@{       |                    �?�O6o3-�?o            `c@������������������������       �                     $@������������������������       ����M��?h             b@~                           �?�G�z��?F             ^@������������������������       �                     "@������������������������       ��Gi����?@            �[@�       �                    �?f���Z�?�           y�@�       �                    �?�{o���?�           P�@�       �                    �?r�q��?�           С@�       �                    �?��.���?I            @\@�       �                     �?���79��?A            @Y@�       �                    �?$��m��?             :@������������������������       �`�Q��?             9@������������������������       �                     �?�       �                    �?��
���?1            �R@������������������������       ���pBI�?/            @R@������������������������       �                      @������������������������       �                     (@�       �                     �?|X&����?V           �@�       �                    �?d"<%�?�           h�@�       �                    �?��W[@k�?�           �@�       �                    �?�lC���?�            �q@������������������������       �$+ޠ�5�?@            @Z@������������������������       �����?u             f@�       �                    �?��4sր�?           pz@������������������������       �        
             2@������������������������       � �[gЯ?�            Py@�       �                    �?��LY�?�            �y@�       �                    �?p^H�&m�?Z            �`@������������������������       ����X�K�?!            �F@������������������������       �        9            @V@�       �                    �?x�>Yd�?�            0q@������������������������       �                      @������������������������       �|)����?�            q@�       �                    �?�:���?�           t�@�       �                    �?�`Y��?x            �f@�       �                    �?6�;�vv�?^            @b@������������������������       �H}m�y��?\            �a@������������������������       �                     @�       �                    �?      �?             B@������������������������       �     ��?             @@������������������������       �                     @�       �                    �?��w��k�?$           8�@�       �                    �?��Nx��?m           P�@������������������������       ���'�`�?k            �d@������������������������       ��d�g��?           @z@�       �                    �?��S�ۿ?�            �q@������������������������       �        -            @R@������������������������       ��|1)��?�            �j@�       �                    �?��>4�g�?            |@�       �                    �?�ݜ�?            �C@�       �                     �?�חF�P�?             ?@������������������������       ������H�?             2@������������������������       ��θ�?             *@������������������������       �                      @�       �                    �?�)���?�            �y@�       �                     �?�%/�A�?�            pp@������������������������       ��2�R�?O            @^@������������������������       ���W3�?Y            �a@�       �                     �?�+�����?W            @b@������������������������       ����"͏�?.            �R@������������������������       �P��E��?)             R@�       �                     �?ܩ���G�?>           ��@�       �                    �?�:�<}=�?�           ��@�       �                    �?�6
����?�           �@�       �                    �?�8��8��?�            �l@������������������������       �ؗp�'ʸ?�            �h@�       �                    �?     ��?             @@������������������������       �r�q��?             @������������������������       �8�Z$���?             :@�       �                    �?��.��?a           Ȁ@�       �                    �?��j�o�?           �y@������������������������       �hA� �?_            �a@������������������������       ��t����?�             q@������������������������       �P�B�y��?T            @_@�       �                    �?ܱ#_��?�            `r@�       �                    �?�t����?            �I@������������������������       �r�q��?             B@�       �                    �?���Q��?             .@������������������������       �                     "@������������������������       �                     @�       �                    �?d�:X�?�            `n@�       �                    �?��p\�?~            �i@������������������������       ��O4R���?             �J@������������������������       �@݈g>h�?^             c@������������������������       �P����?             C@�       �                    �?,����?�           ��@�       �                    �?����j[�?�            �@�       �                    �?4ͧ*���?           h�@������������������������       ��D��S��?.           @}@������������������������       �0 �����?Q            @^@�       �                    �?J�8���?4            �U@������������������������       �z�G�z�?            �A@������������������������       � ��WV�?             J@�       �                    �? ;����?�           P�@�       �                    �?�N,0sm�??           �@�       �                    �?      �?             8@������������������������       �X�Cc�?             ,@������������������������       �ףp=
�?             $@�       �                    �?����Og�?1           �~@������������������������       ���0{9�?�            �t@������������������������       ��Zl�i��?b            @d@�       �                    �?�E����?�            pp@�       �                    �?��H.��?|             i@������������������������       ��(\����?             D@������������������������       ��z�Ga�?g             d@�       �                    �?�G��l��?'            �O@������������������������       �      �?              @������������������������       ��eP*L��?"            �K@�       !                   �?x�s�<��?�           ��@�                          �?hlS���?�	           ��@�       �                    �?���?x.�?�            �@�       �                    �?�!�{QA�?�           ��@������������������������       �                     *@�       �                    �?�c��S��?�           @�@�       �                     �?���?4           �~@�       �                    �?FzW���?�            `r@������������������������       ���|Io��?Q            �]@������������������������       �@�k$��?d            �e@�       �                    �?*S%��?            �h@������������������������       �        9             W@������������������������       �X�Emq�?F            �Z@�       �                    �?���Xh�?�            �k@�       �                     �? ����?-            @P@������������������������       �                     B@������������������������       �XB���?             =@�       �                     �?h�����?c            `c@������������������������       �DrfuN�?<            �W@������������������������       ���7��?'            �N@�       �                    �?P����?�           ̒@������������������������       �                     @�                           �?��ѓ��?�           ��@�                           �?p�Y��?�           ��@������������������������       �8��8��?�             x@������������������������       ��ѯXjy�?�            @s@                         �?8q��^�?)           �@������������������������       �^�!~X�?�            �s@������������������������       ��B!A�?p            �g@                         �?�mA�?Z           ��@                         �?@ѽ�֞?�           p�@������������������������       �        9            �V@                          �?���m�ա?o           ��@	      
                   �?0���|�?�             l@������������������������       �0\�����?w            @f@������������������������       �`Ql�R�?            �G@                         �?���͡?�            0u@������������������������       � M��~?�             q@������������������������       �t�e�í�?'            �P@                          �?to7����?�           $�@                         �?8�����?�           ��@                         �?�P�����?l             e@������������������������       �r�i�+$�?E             [@������������������������       ���Q��?'             N@                         �?����Ԅ�?F           �~@                         �?�������?�             w@������������������������       �                     @������������������������       ���f���?�            �v@������������������������       ��7���?Y             _@                         �?��zi��?            ��@������������������������       �                     @                         �?|뽬��?�           h�@                         �?�q�q�?�             k@������������������������       ��K£���?k             e@������������������������       �"Ae���?            �G@                          �?��v��?r           ��@������������������������       �L�k�)�?           �{@������������������������       �� ���?`            @c@"      +                   �? Լm���?�           û@#      *                   �?�lZ��#}?�           ��@$      '                   �?@v�����?�            �@%      &                    �?�k~X��?�             r@������������������������       �        \            `a@������������������������       � �ޫ��?f            �b@(      )                    �?��a�zt?           ��@������������������������       � �ԍ�m?k           ��@������������������������       ��q�k��v?�           ��@������������������������       �        �            t@,      ;                   �?��8��?            �@-      4                   �?�Ӿjq!�?�           ��@.      1                    �?�����?�           Ѓ@/      0                   �?���؇>�?�            @p@������������������������       �8�B�q�?A            �W@������������������������       �r٣����?d            �d@2      3                   �?��;���?�            `w@������������������������       ���%3�?C            @Y@������������������������       �&>!�q�?�            q@5      8                   �?`�����?S            �@6      7                    �?ཕvt�?@           ��@������������������������       �h4AO+�?%           �|@������������������������       �He��+��?           �z@9      :                    �?05D�b7�?           �@������������������������       ��	]�h��?           �@������������������������       ���k�E��?�           �@<      C                   �?Ї	{�k�?=            �@=      @                    �?n��K�?�            `i@>      ?                   �?�~8�e�?J            �Y@������������������������       ��m����?/            �M@������������������������       �8�$�>�?            �E@A      B                   �?zP1�?K            @Y@������������������������       ���[�p�?#            �G@������������������������       �J��D��?(             K@D      G                    �?pm�n��?�           ��@E      F                   �?�`D��q�?1           0~@������������������������       �     ��?�             p@������������������������       ��C&�l��?�            `l@H      I                   �?�E�%��?w           Ђ@������������������������       ���sK�z�?�            �n@������������������������       �H鮜޹?�            @v@K      �                   �?�q��R�?Q          �A�@L      s                   �?��͉,��?�           ��@M      Z                   �?h%!�!a�?�            �@N      Y                   �?8l�9���?y            �j@O      X                   �?"�
d|�?n            �h@P      U                    �?dWp,���?a            @f@Q      T                   �?�p�o�?�?;            �[@R      S                   �?      �?              P@������������������������       �                     �?������������������������       ����N8�?            �O@������������������������       �"Ae���?            �G@V      W                   �?�萻/#�?&            �P@������������������������       ��\��N��?             C@������������������������       ��c�Α�?             =@������������������������       �                     3@������������������������       �                     1@[      h                    �?DᲯ2�?�           ȕ@\      c                   �?�yD�^�?           P�@]      ^                   �?�*v��??           P~@������������������������       �                     @_      b                   �?{*�?�?<            ~@`      a                   �?�nF$m��?           Pz@������������������������       ���ꤘ�?h             c@������������������������       ���	��j�?�            �p@������������������������       �`��:�?'            �N@d      g                   �?tq�l��?�            Pt@e      f                   �?�-@�w��?�            0p@������������������������       � qP��B�?/            �U@������������������������       ����y�?u            �e@������������������������       �:ɨ��?*            �P@i      p                   �?�ucR�?u           @�@j      m                   �?�yo��4�?%           �|@k      l                   �?@m����?Z            �b@������������������������       �@�E�x�?;            �X@������������������������       �                    �I@n      o                   �?�S_/�m�?�            �s@������������������������       ��-m7"C�?�            �h@������������������������       �x�}b~|�?B            �\@q      r                   �?����5�?P            �^@������������������������       �z�G�z�?$            �K@������������������������       �Pa�.l�?,            �P@t                          �?�*�S���?�           D�@u      |                   �?<��F=]�?y           ��@v      y                   �?f�B���?�            �i@w      x                   �?hx<?v��?K            �]@������������������������       �8�Z$���?            �C@������������������������       �        4             T@z      {                   �?j���� �?9            @U@������������������������       �l��
I��?             ;@������������������������       ���o	��?"             M@}      ~                   �?0��_��?�            0w@������������������������       �`	�<��?e            �a@������������������������       ����^���?�            �l@�      �                   �?�E��&J�?z           ��@�      �                   �?��W���?v             g@�      �                   �?d}h���?.            �Q@������������������������       ������H�?             B@������������������������       ��!���?             A@�      �                   �?���5��?H            �\@������������������������       �      �?$             P@������������������������       �z�G�z�?$             I@�      �                   �?P�cZY�?           �y@�      �                   �? ������?P            �_@������������������������       �                      @������������������������       �0�z��?�?O             _@������������������������       �����,��?�            �q@�      �                   �?Dp{��?c           ��@�      �                    �?�G�
+#�?�           �@�      �                   �?�jTx��?�           P�@�      �                   �?|ܑ��b�?�            pt@�      �                   �?��C���?;            �W@�      �                   �?�㙢�c�?             G@������������������������       �                     @������������������������       ���s����?             E@������������������������       �                     H@�      �                   �?h�1F:�?�             m@�      �                   �?b�2�tk�?             2@������������������������       ��z�G��?             $@������������������������       �                      @�      �                   �?Dw�&��?�            �j@������������������������       �P��BNֱ?f            �d@������������������������       ������?            �H@�      �                   �?���}<S�?0           0~@������������������������       �                     (@�      �                   �?�f���?)           p}@�      �                   �?8��8���?{             h@������������������������       �Xsj�]�?K            @^@������������������������       ���U��?0            �Q@������������������������       �}�rg�?�            pq@�      �                   �?�q�q�?�           `�@������������������������       �        #             J@�      �                   �?V���l�?�           ��@�      �                   �?�_���?v           �@�      �                   �?�ko{޲�?�            �q@�      �                   �?     ^�?K             `@������������������������       ����;QU�?(            @R@������������������������       ��C��2(�?#            �K@������������������������       �`<)�+�?d            @c@�      �                   �?��|�5��?�            �t@�      �                   �?`�I��g�?�            �l@������������������������       �                     @������������������������       ��H�@=��?�            �k@������������������������       ����o_�??             Y@�      �                   �?*X����?K           �@�      �                   �?n�tl��?A            �Z@������������������������       �                     @������������������������       �؁sF���?:             Y@������������������������       �������?
           `y@�      �                   �? �ޚ���?�           �@�      �                    �? F#q��?�           ��@�      �                   �?�S���?           0|@�      �                   �?�X����?V            �`@������������������������       ��}�+r��?;            �W@������������������������       �                    �B@�      �                   �?�@��<�?�            �s@�      �                   �?\-��p�?             =@������������������������       �                     @������������������������       � ��WV�?             :@�      �                   �?P��ʹ�?�             r@������������������������       ���H���?x             h@������������������������       ��9:�l'�?8            @X@�      �                   �?���X��?�            �@�      �                   �?"pc�
�?�            �r@������������������������       �o�U��?�             o@������������������������       �@��8��?"             H@�      �                   �?��
��X�?�            pw@�      �                   �?�ŇG+��?�            �o@������������������������       �r�q��?             @������������������������       ���1��?�            �n@�      �                   �?��}��?M            �^@������������������������       ��#-���?            �A@������������������������       �8�A�0��?8             V@�      �                    �?H'�J7��?�	           
�@�      �                   �?�V8z�	�?[           ,�@������������������������       �@4�1b�?%           0|@�      �                   �?�G:E��?6           @�@������������������������       ����w��?[            �a@������������������������       �Hm6$���?�           ؇@�      �                   �? iS�d�?Y           t�@������������������������       ���swɃ?�           �@�      �                   �?\��m���?�           И@������������������������       ��vΥ�?x            @i@������������������������       ���$���?T           ��@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B�       ��@     ��@    ���@     �@     ��@     .�@    ��@     �@     Ѐ@     0~@     Ѐ@     ~@     ��@     ~@     �{@     @t@      o@     �l@     `h@     @W@     �V@     �c@      @                       @    ���@     x�@    ���@     x�@    ���@     �q@     H�@     �Y@     ��@     @T@     X�@     �@@     @e@      @      R@      @     �X@             �@      =@     �@      7@     ��@      @     �@      H@     �J@      @      0@      @     �B@             p�@     �E@     �k@      @@     ��@      &@     �@      5@     4�@      (@     �N@             @�@      (@     �q@      (@     ؒ@             `�@      "@      5@      �?      @      �?      1@             ��@       @     �Y@      @      @      �?     ʭ@     �f@     j�@      ]@     ��@     �P@      @             ��@     �P@      4@      @     D�@     �O@     ,�@      I@      @@             ��@      I@      @             ��@      I@     ��@     @P@       @             ��@     @P@     �B@             $�@     @P@     x�@      >@     Ѓ@     �A@     p�@     @s@     �y@      e@      @      3@      @      ,@       @      @     �y@     �b@      m@     �T@     �e@     �P@       @             �e@     �P@      q@     �a@       @      (@      �?      "@      �?      @     �p@      `@     `d@     �U@     �Z@     �D@     (�@     x�@     �@     �m@     Й@     �`@     �h@      I@     �f@     �H@     �[@     �A@     �Q@      ,@      0@      �?      "@      �?      @             ��@     �T@     p�@       @      u@      @     �o@      @     �@     �R@      |@     �B@     z@     �B@     @�@      Z@     @@     �O@     t@      G@     �M@     �B@     `p@      "@     `f@      1@      4@      .@     �c@       @     ��@     �D@     0s@      1@      0@      �?     0r@      0@      m@      8@      @             @l@      8@      y@     0r@     �m@     @f@      @      3@      �?      "@       @      $@     `m@     �c@     �`@     @X@     @Y@      O@     @d@     @\@      X@     �M@              $@      X@     �H@     �P@      K@              "@     �P@     �F@     F�@     X�@     ��@     P�@     ��@     �w@      7@     �V@      &@     �V@      "@      1@       @      1@      �?               @     @R@       @     �Q@               @      (@             T�@      r@     ��@     �^@     X�@     �U@      j@     @R@     �B@      Q@     �e@      @     �y@      *@      2@             �x@      *@     @w@     �B@     @^@      *@      @@      *@     @V@             `o@      8@       @              o@      8@     ��@     �d@     �R@     �Z@     �L@     @V@     �J@     @V@      @              2@      2@      ,@      2@      @             X�@      N@     �@     �D@     �d@       @     �w@     �C@     �p@      3@     @R@              h@      3@      q@     �e@      @      A@      @      :@       @      0@      @      $@               @     �p@     �a@     @e@     @W@     �S@     �E@      W@      I@     �X@     �G@      L@      2@     �E@      =@     ��@     ��@     h�@     `w@     p|@     `s@      3@      j@      $@     @g@      "@      7@      @      �?      @      6@     @{@     @Y@     `w@      C@     �`@      @      n@      @@      O@     �O@     �l@      P@      .@      B@      @      >@      "@      @      "@                      @     �j@      <@     �g@      .@      J@      �?     @a@      ,@      9@      *@     ��@     ��@      g@     �~@     �_@     �|@      ,@     `|@     @\@       @     �L@      >@      @      <@      I@       @      �@     @i@     �{@     �Q@      2@      @      "@      @      "@      �?     �z@     @P@     �q@     �H@     @b@      0@     �`@     ``@     �X@     @Y@      �?     �C@     �X@      O@     �@@      >@      @      @      >@      9@     ��@    ���@     ��@     T�@     @s@     P�@     �e@     @�@              *@     �e@     ؀@      ^@     @w@     �R@     �k@      $@     @[@      P@     �[@      G@      c@              W@      G@      N@     �J@     �d@      �?      P@              B@      �?      <@      J@     �Y@      =@     @P@      7@      C@     �`@     ��@              @     �`@     ��@      S@     @�@     �H@     �t@      ;@     �q@     �M@     �{@      E@     @q@      1@     `e@     p@     X�@      $@      �@             �V@      $@     P�@      @     �k@      @     �e@      �?      G@      @     �t@      �?     �p@      @      O@     �n@     H�@     �Y@     x�@      I@     �]@      =@     �S@      5@     �C@     �J@     �{@      E@     �t@              @      E@     Pt@      &@     @\@      b@     �@              @      b@     �@     �V@     �_@     �R@     �W@      0@      ?@      K@     ��@      >@     �y@      8@     @`@     �~@     չ@       @     r�@       @     ��@      @     �q@             `a@      @      b@      @     p�@      �?     ��@      @     ��@             t@     `~@     �@     `u@     H�@     �f@     `|@     �P@     @h@      :@     @Q@      D@     @_@     �\@     @p@      =@      R@     @U@     �g@     @d@     ��@      E@     ��@      5@     �{@      5@     �y@      ^@     (�@      M@     8�@      O@     �@      b@     ��@     �Q@     �`@      F@      M@      =@      >@      .@      <@      ;@     �R@      $@     �B@      1@     �B@     @R@     ��@      D@     �{@      7@      m@      1@     @j@     �@@     ȁ@      ,@      m@      3@     u@     ʧ@     ��@     p�@     ��@     ��@     �l@     �[@     �Y@     �[@     �U@      W@     �U@      P@     �G@      H@      0@              �?      H@      .@      0@      ?@      <@     �C@      4@      2@       @      5@      3@                      1@     ̓@     �_@     `�@      O@     p|@      >@      @             @|@      >@     0y@      2@      c@      �?     `o@      1@     �H@      (@     Pr@      @@     �n@      (@      U@       @     `d@      $@      G@      4@     8�@     @P@     P{@      9@     `b@       @      X@       @     �I@              r@      7@     @g@      *@      Z@      $@     �T@      D@      F@      &@      C@      =@     �^@     \�@      S@     0@     �D@     `d@      @     @\@      @     �@@              T@     �A@      I@       @      3@      ;@      ?@     �A@      u@      3@     �^@      0@     �j@      G@      �@      =@     `c@      .@     �K@      @      @@      &@      7@      ,@      Y@      @      N@      $@      D@      1@     �x@       @      _@               @       @     �^@      .@     �p@     $�@     ��@     ��@     (�@      s@     �@     `p@     @P@      L@      C@       @      C@              @       @      A@      H@             �i@      ;@      @      &@      @      @               @     �h@      0@      d@      @     �C@      $@      E@     �{@              (@      E@     �z@      <@     �d@      @     @]@      8@     �G@      ,@     �p@     �x@     ��@              J@     �x@     ��@     �s@     �r@     �N@     �k@     �K@     @R@      @      Q@      I@      @      @     �b@     �o@     @S@      j@      4@      @             @i@      4@     �E@     �L@     �S@      {@     �M@      H@              @     �M@     �D@      4@      x@     ��@     ��@     h�@     `@     `r@     �c@      E@     �V@      @     �V@     �B@             �o@     �P@      @      9@      @              �?      9@      o@      E@     �e@      3@     �R@      7@     pt@     �u@      K@     `n@      @     @n@     �G@      �?     q@     �Y@     @k@      A@      @      �?     �j@     �@@     �K@      Q@      @      @@      J@      B@     �l@     B�@     �V@     ��@       @     |@     @V@     x�@      M@     �T@      ?@     ��@      a@     b�@      @     �@     �`@     ��@      L@     @b@      S@     x�@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�BHl         �                    �?D���?�e           �@       �                    �?�_q���?|5          �#�@       h                    �?e�(<��?�#           5�@       !                    �?������?�          �@�@                           �?6+3����?P           ��@                           �?��;?Ei�?            D�@       
                     �?L�vD��?w           �@       	                     �?������?�           0�@������������������������       �"��;1Z�?/           P~@������������������������       ���V�-�?�            r@������������������������       ��q�q�?�            �o@                            �?�L#���?�            �p@                           �?��F�D�?z            �h@                           �?@�E�x�?x            �h@                           �?�a�O�?w            @h@������������������������       �����D��?<            @W@������������������������       �        ;            @Y@������������������������       �                      @������������������������       �                      @                           �?b�h�d.�?/            �Q@                           �?`Jj��?(             O@                           �?      �?             @@������������������������       ���� ��?             ?@������������������������       �                     �?������������������������       �                     >@������������������������       �                      @                           �?p��@���?0            @U@                           �? 7���B�?-            @T@������������������������       �        +            �S@������������������������       �                     @                            �?      �?             @������������������������       �                     @������������������������       �                     �?"       Q                    �?8��/ٟ�?J          ���@#       $                    �?H�M�V.�?�          ���@������������������������       �                     @%       B                    �?�}pvc0�?�          ���@&       5                    �? �ߖJ`�?�           �@'       .                    �?$)�U4��?%           ��@(       +                    �?���5��?�           H�@)       *                     �?0�v���?�           ��@������������������������       ��i>���?Z           ��@������������������������       ����]k�?�             l@,       -                     �?p�q��?�             x@������������������������       ��ת2�%�?�            `q@������������������������       �0��_��?D            �Z@/       2                     �?���.�6�?<             W@0       1                    �?�C��2(�?&            �K@������������������������       ��+$�jP�?             ;@������������������������       �                     <@3       4                    �?�?�|�?            �B@������������������������       �P���Q�?             4@������������������������       �        	             1@6       ;                    �?0k�7���?�           H�@7       :                    �?���kx?%	           ��@8       9                     �?��3���?�           X�@������������������������       ��E$���~?X           ��@������������������������       �`a�����?�           x�@������������������������       �        @           $�@<       ?                    �?�X�+Y��?�	           ҭ@=       >                     �?��`qM|�?�           ��@������������������������       ������?�           đ@������������������������       �@U�Sˬ�?�           ��@@       A                     �?P8"y��?�           �@������������������������       �pb@���?R           `�@������������������������       ��yr�?c�?�           x�@C       J                     �?~�HQ��?�           ؇@D       G                    �?PB�~�?           `z@E       F                    �?���.�6�?v             g@������������������������       �HP�s��?]            �b@������������������������       �                     A@H       I                    �?ҳ�wY;�?�            �m@������������������������       ��D�~X�?a             b@������������������������       ����@M^�?:            @W@K       N                    �?�<dVo�?�            Pu@L       M                    �?<�A+K&�?�            �l@������������������������       ����U�?<            �\@������������������������       ����;�?E            �\@O       P                    �?�*�Lk�?J            @\@������������������������       �@-�_ .�?            �B@������������������������       �&:~�Q�?-             S@R       a                    �?�-r~ۓ�?x           0�@S       Z                     �?�ʑ*`�?           ��@T       W                    �?��݉"�?8           �@U       V                    �?�����η?�             l@������������������������       �z�G�z�?             I@������������������������       ���즟E�?j            �e@X       Y                    �? >�֕�?�            �q@������������������������       �                     &@������������������������       ��)2e��?�            �p@[       ^                    �?����?�            �u@\       ]                    �?��0{9�?]            �a@������������������������       ��q�q�?             H@������������������������       ��L��ȕ?A            @W@_       `                    �?�n����?�            �i@������������������������       �                     @������������������������       ��G� �?�            @i@b       e                     �?Z�E����?`             b@c       d                    �?     ��?-             P@������������������������       ����y4F�?             C@������������������������       ��n_Y�K�?             :@f       g                    �?�<ݚ�?3            @T@������������������������       �`���i��?             F@������������������������       ���%��?            �B@i       z                     �?RoQ0�q�?F           ң@j       u                    �?��^�a!�?�           �@k       p                    �?��!�0�?�           ��@l       o                    �?�J�4�?             9@m       n                    �?z�G�z�?             4@������������������������       ��t����?
             1@������������������������       ��q�q�?             @������������������������       �                     @q       r                    �?0�6�0�?�           Ȃ@������������������������       �����>�?�            �r@s       t                    �?v5=�k��?�            s@������������������������       ���8�ͻ�?�             o@������������������������       ��MWl��?&            �L@v       y                    �?�o�8���?           ��@w       x                    �?dAyS��?�           �@������������������������       �0��m0�?            py@������������������������       ��+I�9��?�            �p@������������������������       �D��2(�?p             f@{       �                    �?������?�           ��@|       �                    �?]u�?           x�@}       ~                    �?�m�>���?J           @�@������������������������       �                     �?       �                    �?�����?I           8�@�       �                    �?��0u���?�             n@������������������������       ������H�?             "@������������������������       �h/��y��?�            �l@������������������������       ��sp�1E�?�            ps@�       �                    �?(�-~ ��?�            pt@�       �                    �?`�Q��?^            �b@������������������������       �      �?             @������������������������       �X~�pX��?\            @b@������������������������       ��j��b�?m             f@�       �                    �?����?|            �f@�       �                    �?     ��?*             P@������������������������       �                     @������������������������       ���mo*�?'            �M@������������������������       �Xc!J�ƴ?R            �]@�       �                    �?vϷ���?�           $�@�       �                     �?�����b�?           ��@�       �                    �?�6S-Ņ�?           ��@�       �                    �?�p��f>�?�           ̞@�       �                    �?^Q<��K�?3           P�@�       �                    �?H�3��q�?�           �@�       �                    �?�<ݚ�?b             c@������������������������       ��<ݚ�?\             b@������������������������       ��<ݚ�?             "@�       �                    �?(�?P��?(           `�@������������������������       ��i�,�;�?�             x@������������������������       ���<D�m�?8           �~@�       �                    �?��Lu-��?�            �p@������������������������       ���z*�o�?b            �c@������������������������       �Dc}h���?G             \@�       �                    �?�7�^�?�           ��@�       �                    �?n��K�?{            `i@������������������������       ����!pc�?             &@������������������������       �     8�?u             h@������������������������       �ȑ����?2           @}@�       �                    �?J�땐��?3           x�@�       �                    �?�fq
B.�?Q           ��@�       �                    �?@@c�w�?�           ��@�       �                    �?�Q��k�?3             T@������������������������       �z��R[�?.            �Q@������������������������       �                     $@�       �                    �?p�_����?�            �@������������������������       ���6���?�            p@������������������������       �X�?�ݾ?           0z@�       �                    �?�҇���?k            �g@������������������������       �      �?             (@������������������������       �HN�z��?d             f@�       �                    �?���!�?�            �v@������������������������       � pƵHP�?%             J@�       �                    �?4O��n�?�            �s@������������������������       �      �?'             Q@������������������������       �����X��?�            �n@�       �                    �?d��x��?            ^�@�       �                    �?R���6�?�           @�@�       �                    �?�Je\���?f            @d@�       �                    �?4�M�f��?B            �Y@�       �                    �?�q�q��?>             X@�       �                    �?��.k���?8            @U@������������������������       �      �?              @������������������������       ���}E��?6            �T@������������������������       �"pc�
�?             &@������������������������       �                     @�       �                    �?�G�z��?$             N@�       �                    �?�w��#��?             I@������������������������       ��lg����?            �E@������������������������       �؇���X�?             @������������������������       �                     $@�       �                    �?��!Y��?           ��@�       �                    �?�+��<v�?�           ȇ@�       �                    �?��m����?z           ��@������������������������       �`=��?��?�            �p@������������������������       � ��&*6�?�            0t@������������������������       �r�᮹��?b             e@�       �                    �?� �i��?@           P@�       �                    �?8��H��?            y@������������������������       ������?[             a@������������������������       ��U�=���?�            �p@������������������������       �Fn�圴�?<            @Y@�       �                    �?�S	���?~           |�@�       �                    �?��8����?�           ��@������������������������       � h'M#�?e            �f@�       �                    �?0�A�A��?N           ؀@������������������������       ��^�����?7            �U@������������������������       �ps�r��?           P|@�       �                    �?�H�@=��?�            �t@������������������������       �                     F@�       �                    �?�����?�            r@������������������������       ��r����?            �F@������������������������       �\#r��?�            �n@�       �                    �?��q�m�?�           ��@�       �                    �?��>���?�           �@�       �                    �?�?�'�@�?-           �|@�       �                    �?B� ��?-            �Q@�       �                     �?�-ῃ�?(            �N@������������������������       ���S���?             >@������������������������       ��n`���?             ?@������������������������       �                     "@�       �                    �?��h�V�?             x@�       �                     �?�Μ�5�?M            �[@������������������������       ����U�?+            �L@������������������������       �        "             K@�       �                     �?�4�)w�?�            0q@������������������������       �x�}b~|�?q            `e@������������������������       � ��WV�?B             Z@�       �                     �?�F~���?m            �f@�       �                    �?��6���?6             U@������������������������       �                     @������������������������       ����;+"�?4            �S@�       �                    �?D]��;��?7            @X@������������������������       �                     "@������������������������       �d�
��?0             V@�       �                    �?`���pR�?�           8�@�       �                     �?�h����?e             e@������������������������       �@uvI��?:            �X@������������������������       ���?^�k�?+            �Q@�       �                    �?�����H�?�           ��@�       �                     �?
�c�Z�?B             Y@������������������������       ����Q��?"            �K@������������������������       ����V��?             �F@�       �                     �?�S(��d�?H           ؀@������������������������       � �_�x�?�            `o@������������������������       ��n���?�             r@�       �                   �?tK�r_��?0          ��@�       O                    �?��ӣ��?�          ���@�       4                   �?X�����?}           -�@�                          �?�{�/���?p           ��@�                          �?��O5���?_           p�@�                          �?�P�*�?�           X�@�                          �?�m�!�?�            �r@                          �?��>4և�?K             \@������������������������       �l��
I��?             ;@������������������������       ��ģ�a@�?;            @U@                         �? ������?{            �g@������������������������       �                     @������������������������       ��x�V�?x             g@                         �?��8�<�?�            �u@������������������������       �ܑ-Z���?�            �j@������������������������       � =[y��?W             a@	                         �?b �57�?�           ��@
                         �? 7���B�?             ;@������������������������       �                     0@������������������������       ��C��2(�?             &@                         �?���>{�?�           ��@������������������������       ���h�V�?�             x@������������������������       ��ѯXjy�?�            @s@      #                   �?�v�g1��?           ��@                         �?v�_���?�            �m@                         �?��qC�?0            �S@                         �?��0{9�?            �G@������������������������       �                     �?                         �?*
;&���?             G@������������������������       ��T|n�q�?            �E@������������������������       �                     @                         �?     ��?             @@������������������������       �l��
I��?             ;@������������������������       �                     @                          �?��t���?c            �c@                         �?0�й���?Z            @b@                         �?���y4F�?             C@������������������������       �                     @������������������������       �      �?             @@������������������������       �h�WH��?B             [@!      "                   �?r�q��?	             (@������������������������       �      �?              @������������������������       �                     @$      -                   �?��b�h8�?~           ��@%      &                   �?�.ߴ#�?^           (�@������������������������       �                     @'      *                   �?x/ ��?[           �@(      )                   �?��Y�\ܻ?�            �t@������������������������       �        7            @T@������������������������       �x���<�?�             o@+      ,                   �?�&�� .�?�             k@������������������������       �        !            �K@������������������������       �H�!b	�?g            @d@.      1                   �?,4k@���?            0}@/      0                   �?�IєX�?~            �i@������������������������       �        #             O@������������������������       �@�j;��?[            �a@2      3                   �?�?�(|�?�            pp@������������������������       �`2U0*��?!             I@������������������������       �(�݂��?�            �j@5      >                   �?��-�=��?           ��@6      ;                   �?��R�?z           Ȏ@7      :                   �?@ԕ���?�           �@8      9                   �?��کd�?�            �i@������������������������       �                     ;@������������������������       ��Y�ߠ?u            `f@������������������������       ��f�Ibp?D           0@<      =                   �?��Q���?�            �q@������������������������       �䯦s#�?H            �Z@������������������������       ��s��9n�?j            �e@?      F                   �?H���C`�?�           L�@@      C                   �?L]n�!�?�             n@A      B                   �?�Ŗ�Pw�?^            @a@������������������������       �����?�?            �F@������������������������       �        B            @W@D      E                   �?x�K��??            �Y@������������������������       ��n_Y�K�?"             J@������������������������       ����Q��?             I@G      L                   �?����{�?�           �@H      K                   �?�Ę�;�?x            �g@I      J                   �?@�n���?E            �Y@������������������������       �                     "@������������������������       ���K2��??            �W@������������������������       ����!pc�?3             V@M      N                   �?�z�r��?~            �@������������������������       � dϛ�p?*           @~@������������������������       �     ��?T             `@P      �                   �?d�K�[��?)           b�@Q      l                   �?��Ց��?           ��@R      _                   �?Шݛ��?�           �@S      ^                   �?p�^����?�            �w@T      [                   �?�f�l$�?�            �v@U      X                   �?�U���?�            �o@V      W                   �?�Ń��̧?4             U@������������������������       ��(\����?2             T@������������������������       �                     @Y      Z                   �?ҳ�wY;�?n            @e@������������������������       �4�B��?[            �b@������������������������       ��eP*L��?             6@\      ]                   �?���>4ֵ?=             \@������������������������       �                     =@������������������������       � ,U,?��?,            �T@������������������������       �        	             0@`      a                   �?`xA�X�?�            �@������������������������       �                     @b      g                   �?8i�w1l�?�           �@c      f                   �?��s}n�?�            �t@d      e                   �?��.��C�?�             q@������������������������       �����?s             f@������������������������       ���8�$>�?;            @X@������������������������       �,�+�C�?"            �K@h      i                   �?�c:��?�           ��@������������������������       � �ZH���?�            0y@j      k                   �?�IєX�?           �z@������������������������       �P��a4�?y            �g@������������������������       � 1�/Gu�?�            �m@m      x                   �?&�����?Q           @�@n      q                   �?��r2�M�?g           Ў@o      p                   �?@N�4��?r           ��@������������������������       ��ۏ��?'           �~@������������������������       � >�֕�?K            @Z@r      u                   �?|�y]%��?�            �x@s      t                   �? V�����?�            �r@������������������������       �^H���+�?            �B@������������������������       �`��F:u�?�            Pp@v      w                   �?��s��?8            �W@������������������������       ��7��?            �C@������������������������       �h�����?!             L@y      ~                   �?<�Q��P�?�           ��@z      }                   �?4�2%ޑ�?            �A@{      |                   �?�E��ӭ�?             2@������������������������       ��z�G��?             $@������������������������       �      �?              @������������������������       �@�0�!��?	             1@      �                   �? ���]�?�           ��@������������������������       �b�����?�             u@�      �                   �?�&��e��?�            x@������������������������       ��ma�H��?c             c@������������������������       �\I���?�?�             m@�      �                   �?|��#���?"	           �@�      �                   �?�%�r��?           ��@�      �                   �?�5?'L{�?�           h�@�      �                   �?�]�h\��?           �z@�      �                   �?0�z��?�?�            @w@������������������������       �        ,            �P@������������������������       ����J��?�             s@�      �                   �?XB���?$             M@������������������������       �                     @������������������������       �h㱪��?#            �K@�      �                   �? Qr�?�           ��@������������������������       � ;гQ�v?�           ��@������������������������       �0�ޤ��?Q            @`@�      �                   �? M���j?           ��@�      �                   �?�������?�            �k@������������������������       �                     C@������������������������       �@t�!�a�?x            �f@������������������������       � ��ɀ�_?�           4�@�      �                   �?H,���?           H�@�      �                   �?l`N���?�            �s@�      �                   �?���?�            `l@������������������������       ��d��Pb�?o            @f@������������������������       ����Q �?!            �H@������������������������       �`Y���?8            �V@�      �                   �?�2>�w0�?K           X�@�      �                   �?6�Ee�?�            �t@������������������������       ��I�b�?�            �p@������������������������       ����Q��?$            @P@������������������������       �P����?}            �g@�      �                   �?�Z����?y           ˾@�      �                   �?P�/��??           ��@�      �                   �?�	O��?H           �@�      �                   �?�z[�<��?           �z@�      �                    �?@-�_ .�?            �B@�      �                   �?���N8�?             5@������������������������       ���S�ۿ?	             .@������������������������       �                     @�      �                   �?      �?             0@������������������������       ��8��8��?	             (@������������������������       �                     @�      �                    �?���Ԥ�?�            �x@�      �                   �?��fq��?z            �g@������������������������       ��LQ�1	�?E            �\@������������������������       ��I�w�"�?5             S@�      �                   �?�g��@(�?�            @i@������������������������       ��	j*D�?]            �a@������������������������       ���Q:��?&            �M@�      �                    �?�LLb��?3           @@�      �                   �?�������?~            `j@�      �                   �?�+$�jP�?             ;@������������������������       ���<b���?             7@������������������������       �                     @�      �                   �?H��	,U�?k             g@������������������������       �L�];�?S            �a@������������������������       �0,Tg��?             E@�      �                   �?.s��J�?�            r@�      �                   �? �Cc}�?!             L@������������������������       �`2U0*��?             I@������������������������       ��q�q�?             @�      �                   �?��^���?�             m@������������������������       ��!d��?r            �f@������������������������       ���.k���?"            �I@�      �                   �?�q�s��?�            Px@�      �                    �?`׀�:M�?-            �R@�      �                   �? 7���B�?             ;@������������������������       �                     $@������������������������       ��IєX�?             1@������������������������       �                    �G@�      �                    �?v�>��?�            �s@�      �                   �?F�E���?_            �a@������������������������       �:	��ʵ�?            �F@������������������������       ��J��%�?@            �X@�      �                   �?�+��<��?k            �e@������������������������       �@�&b
}�?3            �U@������������������������       �:�1�(��?8            @U@�      �                    �?�	1��Ѽ?:           ��@�      �                   �?Х���?�           f�@�      �                   �?ĵtHA��?           ��@�      �                   �?���E0�?�            Px@������������������������       �                     @������������������������       �8��X��?�            �w@������������������������       ��D�ғ�?           ��@�      �                   �?@�&��?�           H�@�      �                   �?�����?�            0x@������������������������       �0��P�?e            �d@������������������������       �(�y�?�            �k@�      �                   �?�=����?�           <�@�      �                   �?�F��O�?�            @r@������������������������       �                     �?������������������������       �DE�SA_�?�            0r@������������������������       �dO6�]�?�           X�@�      �                   �?X�R�m^�?�	           �@�      �                   �?���	�?           $�@�      �                   �?,N�_� �?
           �{@������������������������       �                      @������������������������       ��>	<2�?	           �{@������������������������       ��v��?           4�@�      �                   �?��ǘ}�?�           С@�      �                   �?��|�N
�?>           8�@�      �                   �?2%ޑ��?_            �a@������������������������       �                      @������������������������       �0)RH'�?^            @a@������������������������       �P������?�            �w@�      �                   �?觇Z�1�?`           ��@�      �                   �?��au��?           �{@������������������������       �                     @������������������������       ��d�m븿?           P{@������������������������       ������?\           ��@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B�       k�@     ��@    ���@     ��@     �@     ��@     >�@     �@     @�@     �@     Ȉ@     �@     �@     �~@     �|@     �s@     Pq@      j@     `f@     �[@     @U@     @e@     �o@      0@     @h@      @      h@      @      h@       @     �V@       @     @Y@                       @       @              M@      (@      M@      @      <@      @      ;@      @      �?              >@                       @     �S@      @     �S@      @     �S@                      @      �?      @              @      �?             ��@     �@     ��@     �@      @             ��@     �@     ��@     �p@     X�@      V@      �@     �T@     ��@      N@     ��@      :@     �g@      A@     �v@      6@     �p@      (@      X@      $@     �U@      @      I@      @      6@      @      <@              B@      �?      3@      �?      1@             ��@     �f@     ��@      &@     ,�@      &@     ��@      @     H�@      @     $�@             ��@      e@     (�@      V@     �@      L@     ��@      @@     ؝@     @T@     ē@     �C@     (�@      E@     �d@     ��@      X@     `t@      (@     �e@      (@     @a@              A@      U@     @c@      H@     @X@      B@     �L@      Q@     q@     �C@     �g@      @     �[@     �A@     �S@      =@      U@       @     �A@      ;@     �H@     �@     �d@     ��@     �K@     �}@      ;@     �j@      &@      D@      $@     �e@      �?     �p@      0@      &@             �o@      0@      t@      <@      ^@      5@      <@      4@      W@      �?      i@      @      @             `h@      @      B@     @[@      2@      G@       @      >@      $@      0@      2@     �O@      �?     �E@      1@      4@     p�@     l�@     (�@     ��@     Pz@     �i@      @      5@      @      0@       @      .@       @      �?              @     z@      g@      k@      T@      i@      Z@     �c@     �V@      F@      *@      X@     ��@     @R@     Ȃ@     �E@     �v@      >@     �m@      7@      c@     �x@     ��@     pu@     ��@     �k@     �t@      �?             �k@     �t@     �e@      Q@      �?       @     `e@      N@      I@     Pp@      ^@     �i@     �Y@      H@       @       @      Y@      G@      2@     �c@      I@     �`@     �F@      3@              @     �F@      ,@      @     @\@     �@     F�@     ��@     b�@     $�@      �@     đ@     �@     �@     ps@     ��@     �Q@     �]@      A@      \@      @@      @       @     8�@     �B@     �w@      @     �|@      >@      ?@      n@       @     �c@      =@     �T@     �b@     X�@     �`@     �Q@      @       @      `@     �O@      0@     @|@     ��@     `|@     P�@     �`@     H�@     �E@     �P@      *@     �L@      *@      $@             0�@      >@     �o@      @     �x@      ;@     @X@     �V@      @      @     �V@     @U@      G@      t@      �?     �I@     �F@     �p@      1@     �I@      <@     @k@     �@     ��@     ��@     �l@     �T@      T@     �H@     �J@     �H@     �G@      D@     �F@      �?      �?     �C@      F@      "@       @              @     �@@      ;@     �@@      1@      ;@      0@      @      �?              $@     h�@     �b@     ��@     @W@     H�@     �C@     Pp@       @     @r@      ?@     �\@      K@     �{@     �K@     �w@      7@     �`@      @     �n@      4@     @Q@      @@     �V@     (�@      N@     ��@       @     �f@      M@     ~@      :@      N@      @@     Pz@      >@     �r@              F@      >@     0p@      @     �C@      8@     �k@     ��@     ��@     �~@     �b@     �x@      N@      ?@     �C@      6@     �C@      0@      ,@      @      9@      "@             �v@      5@     @[@       @     �K@       @      K@              p@      3@     �c@      .@      Y@      @      W@     @V@      G@      C@              @      G@     �@@      G@     �I@              "@      G@      E@     �R@     �@      @     �d@      �?     @X@       @      Q@     �Q@     ��@      =@     �Q@      6@     �@@      @      C@      E@     @      6@     �l@      4@     �p@     ��@    ���@     P�@     ?�@     �@     t�@     F�@     ��@     h�@      t@     �w@     q@     �l@     �Q@      F@      Q@       @      3@      B@     �H@     @g@      @      @             �f@      @     �b@     @i@      2@     �h@     @`@      @      �@     �H@      :@      �?      0@              $@      �?     0�@      H@     �v@      5@     �q@      ;@     $�@     �k@     @T@     �c@     �J@      :@      D@      @      �?             �C@      @      B@      @      @              *@      3@       @      3@      @              <@     @`@      2@      `@       @      >@              @       @      8@      $@     �X@      $@       @      @       @      @             ��@      P@     P�@      ;@      @             8�@      ;@     `s@      3@     @T@             �l@      3@      j@       @     �K@             @c@       @     �z@     �B@      h@      (@      O@             @`@      (@     �m@      9@      H@       @     �g@      7@      j@     p�@     @T@     @�@      @     �@      @     `i@              ;@      @      f@      �?      @     @S@     `i@      D@     �P@     �B@      a@     �_@     ��@     �D@     �h@      �?      a@      �?      F@             @W@      D@      O@      4@      @@      4@      >@     �U@     h�@      9@     �d@      �?     �Y@              "@      �?     @W@      8@      P@     �N@     8�@      �?     0~@      N@      Q@     ��@     �@     "�@     �@     <�@     pw@     �T@     �r@     �P@     �r@      O@      h@       @     �T@       @     �S@              @      N@     �[@      H@      Y@      (@      $@      @     �Z@              =@      @     �S@      0@             �@      S@      @             �@      S@     �s@      *@     �p@      "@     �e@      @     @W@      @     �I@      @     �@     �O@     �v@      C@      y@      9@      f@      &@     �k@      ,@     �@     p�@     �m@     p�@      ^@     �}@      5@     0}@     �X@      @      ]@     Pq@      9@     q@      *@      8@      (@      o@     �V@      @     �B@       @      K@       @     ��@      X@      ;@       @      *@      @      @      @      @       @      ,@      @     ؃@      V@     �q@      L@     v@      @@     �a@      *@     �j@      3@     �t@     ��@      0@     f�@      ,@     0�@       @     `z@      @     �v@             �P@      @     �r@       @      L@              @       @     �J@      @     ��@      @     ��@      @     �_@       @     ��@      �?     `k@              C@      �?     �f@      �?     0�@     �s@     h�@     �`@     @g@     �U@     �a@     @Q@     @[@      1@      @@      G@     �F@      g@     0u@     �]@     �j@     @W@     �e@      :@     �C@     @P@     @_@     D�@     z�@     @�@     ��@      �@      z@     �p@     �c@       @     �A@      �?      4@      �?      ,@              @      �?      .@      �?      &@              @     �p@      _@     �`@      M@     �R@      D@      M@      2@      a@     �P@     �X@      F@     �B@      6@      n@     0p@     �]@     @W@      @      6@      @      2@              @     @\@     �Q@     �T@      N@      ?@      &@     �^@     �d@      @      I@       @      H@      @       @     @]@      ]@     @W@     @V@      8@      ;@      i@     �g@      �?     @R@      �?      :@              $@      �?      0@             �G@     �h@      ]@     �Y@      D@     �B@       @     �P@      @@      X@      S@     �H@      C@     �G@      C@     �x@     �@      e@     �@     �W@     �@     �F@     �u@              @     �F@      u@     �H@     X�@     �R@     �@      4@     �v@      $@     @c@      $@     �j@     �K@     ��@      8@     �p@              �?      8@     �p@      ?@     `�@      l@     "�@     �S@     �@      >@     �y@               @      >@     �y@     �H@     p�@      b@     ��@      E@     �}@      6@     �]@               @      6@      ]@      4@     pv@     �Y@     �@      =@     �y@              @      =@     �y@     �R@     |�@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�B�h         
                   �?�
{�(��?He           �@       �                    �?DU���?�4          ���@       "                    �?��E�7�?�#           _�@                           �?���~h�?<           ��@                           �?^��+��?�           T�@                           �?\�ߢG��?�           P�@                           �?�)�8��?�            �@                            �?"��h��?`           �@	       
                     �?̔�&E��?�           ��@������������������������       ��ćo��?           @|@������������������������       �lutee�?�            �p@������������������������       ��'�H��?�            �m@                            �?؀���˲?V            ``@������������������������       �        B            �X@������������������������       �6YE�t�?            �@@                           �?P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                     �?                           �?���'Z��?y            �i@                            �?��I�~R�?u            �h@                           �? �}�$>�?V            �a@                           �?@��8��?:             X@                           �?`Ql�R�?8            �W@������������������������       �        7             W@������������������������       �                      @������������������������       �                      @������������������������       �                    �G@                           �?H�ՠ&��?             K@������������������������       �                    �G@������������������������       �                     @        !                    �?և���X�?             @������������������������       �                     @������������������������       �                     @#       f                    �?��jE��?�           ���@$       C                    �?0��oj�?�          �'�@%       :                    �?�(�d�?�           ��@&       /                     �?`v�FW��?o           ��@'       (                    �?��w�Z�?a           ��@������������������������       �                      @)       .                    �?`�1of�?_           ��@*       -                    �?8�H��?<           p�@+       ,                    �?����Aٴ?"           0�@������������������������       �@ �Z�?i           X�@������������������������       ��u��X�?�            �s@������������������������       �      �?             D@������������������������       �        #            @Q@0       7                    �?���K��?           �z@1       2                    �?Zy'��?�            �x@������������������������       �                     @3       6                    �?�>p��+�?�            px@4       5                    �?`�3Ka��?�            �u@������������������������       �s�pz�?�             n@������������������������       �,�+�C�?G            �[@������������������������       ��G�z��?             D@8       9                    �?�g�y��?             ?@������������������������       �$�q-�?
             *@������������������������       �                     2@;       <                    �?*
;&���?             G@������������������������       �                     9@=       @                    �?�q�q�?             5@>       ?                     �?��
ц��?             *@������������������������       �      �?             @������������������������       �և���X�?             @A       B                     �?      �?              @������������������������       �z�G�z�?             @������������������������       �                     @D       [                    �?�+�'��?I          �Q�@E       P                     �?p}g@{`�?           ���@F       M                    �?�����?�           ֵ@G       J                    �?�~����?�           ��@H       I                    �? y�ݒ�o?l           ��@������������������������       � ��^)~?e           $�@������������������������       �                   В@K       L                    �?HY��Ũ�?           B�@������������������������       �p�B��?�           ��@������������������������       ���pBI�?<           ��@N       O                    �?��W3�?o           ��@������������������������       ��%o��?�            �t@������������������������       ����8���?�             m@Q       X                    �?�;�̿?1           �@R       U                    �?���԰?<           ��@S       T                    �?���°�?�           ��@������������������������       � �#F���?�           h�@������������������������       �        4           �@V       W                    �? >�֕�?{           ��@������������������������       �ȳ�"k�?�           ��@������������������������       �h���Bx�?�           (�@Y       Z                    �?Z.q2�7�?�            @y@������������������������       ��>:���?�            `l@������������������������       �ڵ��~!�?d             f@\       c                    �?���٩d�?)           Њ@]       `                     �?@Z�Ћx�?�           ��@^       _                    �?K�.�?!           �{@������������������������       � ������?s            �g@������������������������       �PYR�?�             p@a       b                    �? �q�q�?�             r@������������������������       �        ;            @V@������������������������       �����9�?�            �h@d       e                     �?���� �?M            �^@������������������������       ��M���?)             Q@������������������������       ���N`.�?$            �K@g       x                     �?���9��?�           ��@h       s                    �?�E�S�?5           �@i       n                    �?8�Z$���?�           x�@j       m                    �?�.k/&��?�           ��@k       l                    �?�輚�?�            Pr@������������������������       ��|K��2�?M             `@������������������������       ���p �?c            �d@������������������������       ��]3m��?�            0y@o       r                    �?��swʭ�?�            `z@p       q                    �?������?U            �c@������������������������       �                     J@������������������������       �^%�e��?<            �Z@������������������������       �@v�禺�?�            �p@t       w                    �?z�G�z�?�            �k@u       v                    �?�ɞ`s�?,            �N@������������������������       ��㙢�c�?             7@������������������������       �\�Uo��?             C@������������������������       �">R��?f            �c@y       �                    �?�N��D�?�           P�@z                           �?�S�w���?�           x�@{       |                    �?�Ԝ7�?H           `�@������������������������       �����w�?D            @[@}       ~                    �?��2��?           �y@������������������������       �z�����?E            �]@������������������������       ���[�?�            �r@�       �                    �?L� P?)�?�            0r@�       �                    �?���Q �??            �X@������������������������       ��:�^���?            �F@������������������������       �X�Emq�?"            �J@������������������������       �(S��C��?v             h@�       �                    �?��^ҺR�?�            �l@������������������������       �`'�J�?            �I@�       �                    �?�(̶h�?k            @f@������������������������       ��<ݚ�?             B@������������������������       �,�d�vK�?U            �a@�       �                    �?&�����?�           Ժ@�       �                    �?��lF��?�           F�@�       �                    �?�/e�U��?           �@�       �                    �?L������?_            @b@�       �                    �?����?K            @\@�       �                    �?��hq��?E            �Z@�       �                     �?ܾ�z�<�?B             Z@������������������������       �      �?             8@������������������������       �x�G�z�?1             T@�       �                     �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                    �@@�       �                     �?f`q�)�?�           ̐@�       �                    �?��Jr���?Q           0�@�       �                    �?��t��?           �|@�       �                    �?�ʻ����?]             a@������������������������       �4�M�f��?C            �Y@������������������������       �H�V�e��?             A@�       �                    �? �)���?�            @t@������������������������       � pƵHP�?v             j@������������������������       �        I             ]@�       �                    �?�z�G��?5            �V@������������������������       �      �?             B@������������������������       �                      K@�       �                    �?�i�c�~�?[           h�@�       �                    �?�+̸�?�            `l@�       �                    �?      �?k             e@������������������������       �U�T��?V             a@������������������������       ����@M^�?             ?@������������������������       �@�r-��?(            �M@�       �                    �? �\���?�            �r@�       �                    �?pU:6Y�?�            p@������������������������       �����?�?u            �f@������������������������       ��g<a�?8            @S@������������������������       ���p\�?            �D@�       �                    �?M����?|           ��@�       �                    �?�q�i�?�            �@�       �                     �?�X���?             F@�       �                    �?r�q��?             8@������������������������       �        	             &@������������������������       �                     *@�       �                    �?z�G�z�?             4@������������������������       �                     @������������������������       ��IєX�?             1@�       �                    �?�e�U�?�           P�@�       �                    �?h�U�_˾?�           H�@������������������������       �                     @�       �                     �?`Jj��?�           0�@������������������������       ��-�[�?�            �x@������������������������       � ,��-�?�            �y@�       �                     �?vH_-�m�?�            �r@������������������������       ��Y�R_�?S            �a@������������������������       �,��c{�?W            �c@�       �                    �?�������?�           x�@�       �                    �?��?
           �@�       �                    �? 7���B�?             ;@������������������������       �                      @�       �                     �?�}�+r��?
             3@������������������������       ������H�?             "@������������������������       �                     $@�       �                    �?�̏�i�?�           �@�       �                     �?�%IM��?           pz@������������������������       ��:�^���?�            @m@������������������������       ����N8�?w            �g@�       �                     �?��A����?�            �w@������������������������       � �r�ѷ?o             g@������������������������       ���S�ۿ?y            `h@�       �                     �?t�z|�?�            r@�       �                    �?��c����?R             a@�       �                    �?�I�w�"�?.             S@������������������������       �                     @������������������������       �tk~X��?,             R@�       �                    �?��7��?$            �N@������������������������       �                      @������������������������       ��#ʆA��?            �J@�       �                    �?:�lO�?b             c@�       �                    �?�û��|�?.            @Q@������������������������       �                     @������������������������       ��q�q�?*            �O@�       �                    �?�L"p�?4            �T@������������������������       �        	             (@������������������������       ���U��?+            �Q@�       �                    �?t�0�k�?R           b�@�       �                    �? �5yy�?a            �@������������������������       �        O            @b@�       �                    �?��V9��?           p�@�       �                     �?�r��Ł?           �|@������������������������       �@�:;��?o            �f@������������������������       ��yf��\}?�            `q@�       �                     �?����Ʃ?�            0x@�       �                    �?�ۊ�̴?e            �d@������������������������       ����.�6�?             G@������������������������       �0x�!���?G            �]@�       �                    �?`׀�:M�?�            �k@������������������������       �@3����?!             K@������������������������       � ��N8�?m             e@�                          �?�@ ��?�           ��@�       �                    �?� ? ��?�           ��@�       �                     �?     x�?�             x@�       �                    �?�w���?d            @d@������������������������       �Dc}h��?E             \@������������������������       ���H�}�?             I@�       �                    �?�As`�?�            �k@������������������������       �t�����?n             e@������������������������       �X�<ݚ�?             K@�       �                    �?�B ���?�           ��@�       �                     �?�I�Aǫ�?
           p�@�       �                    �?��D���?�             x@������������������������       �                      @������������������������       �     ��?�             x@�       �                    �?ଵێ�?           �z@������������������������       �                     @������������������������       ����w�C�?           Pz@�       �                     �?t�U����?�            �t@������������������������       �|�M���?i            @e@�                           �?lGts��?o            �d@������������������������       �                     @������������������������       ������H�?m            @d@                         �?�F����?           ��@������������������������       �                     .@                         �?�p�_�:�?           (�@                          �?�ՙ�?m             e@������������������������       ����|���?0            @S@������������������������       �t]����?=            �V@      	                    �?�\�D��?�           �@������������������������       �     >�?�             p@������������������������       �����˵�?           �y@      �                   �?�QпYt�?�0          �U�@      k                   �?��BZ���?�           H�@      >                   �?�CQ	C�?�           p�@      /                   �?0F��u�?�           .�@                          �?��E�h��?!           ��@                         �?<{����?Y           �@������������������������       �      �?             @                         �?��ճC|�?W            �@                         �?`��qO�?           ��@                          �?�q�q�?�            �o@������������������������       �d,���O�?_             c@������������������������       ���e�B��?=            �Y@                          �?@bC�Ҥ?�           ��@������������������������       � d��F��?�            u@������������������������       ��ъ��h�?�            r@                          �?XC2 ��?;           x�@                         �?��P~/j�?�            �t@������������������������       �">�֕�?-            �Q@������������������������       � ����~?�            �p@                         �?h2��v�?t             h@������������������������       ���.k���?             A@������������������������       �        ^            �c@!      (                    �?�C�i��?�           �@"      %                   �?�������?           p{@#      $                   �?`	<J���?�            Pu@������������������������       ������?�            �i@������������������������       ��\=lf�?T            �`@&      '                   �?d}h���?:            �X@������������������������       �J�8���?             =@������������������������       ���.N"Ҭ?'            @Q@)      ,                   �?�(ȋ'�?�           �@*      +                   �?����?�           `�@������������������������       �P�tj״?1           �~@������������������������       � ,V�ނ�?R            �_@-      .                   �?П[;U��?3            �U@������������������������       ���[�p�?            �G@������������������������       �P���Q�?             D@0      7                   �?��d��?�           Ȅ@1      4                   �?���.��?           �z@2      3                    �?���L��?+            �Q@������������������������       �d��0u��?             >@������������������������       �R���Q�?             D@5      6                    �?p�G�:	�?�            �v@������������������������       � 	��p�?@            �U@������������������������       ����{}̳?�            q@8      ;                   �?�6L"�?�            `m@9      :                    �?��v$���?O            �^@������������������������       ��(\����?3             T@������������������������       �                     E@<      =                    �?���͡?>            @\@������������������������       ��&=�w��?            �J@������������������������       �                     N@?      T                   �?|r��!�?�           ��@@      I                    �?������?�           T�@A      D                   �?��4�w��?�           <�@B      C                   �?8�Z$���?             *@������������������������       ��<ݚ�?             "@������������������������       �                     @E      H                   �?t���Ú�?�           �@F      G                   �?h�z��?2           ��@������������������������       ��>s{Ab�?           `}@������������������������       ��\�D��?           �{@������������������������       ��y��*�?j            �e@J      O                   �?��|�#��?�           0�@K      N                   �?���y4F�?             3@L      M                   �?������?             .@������������������������       ��z�G��?             $@������������������������       �z�G�z�?             @������������������������       �                     @P      Q                   �?�!�'�?�           ��@������������������������       ����2"��?�             x@R      S                   �?@;�"�?�            w@������������������������       �V^���?�            �p@������������������������       �$�q-�??             Z@U      `                    �?l"
{���?r           �@V      [                   �?�)�=���?�           ȃ@W      Z                   �?؇���X�?             5@X      Y                   �?@�0�!��?
             1@������������������������       �"pc�
�?             &@������������������������       �r�q��?             @������������������������       �                     @\      ]                   �?�psy&�?�            �@������������������������       ��/5mvq�?�             s@^      _                   �?�kb97�?�            @s@������������������������       ��&/�E�?W             _@������������������������       � �r�ѷ?v             g@a      f                   �?p���^�?�           X�@b      e                   �?�I�w�"�?             C@c      d                   �?�LQ�1	�?             7@������������������������       ��t����?             1@������������������������       �      �?             @������������������������       ���S�ۿ?	             .@g      h                   �?`u>�)�?�           (�@������������������������       ��9����?�            �t@i      j                   �?�/a��I�?�            �y@������������������������       �@�#����?d             d@������������������������       �0*��ɾ?�             o@l      {                   �?^�m,��?�           `�@m      t                    �?�'t���?�           ȇ@n      q                   �?������?�            �v@o      p                   �?|��?���?�             k@������������������������       �8�Z$���?             *@������������������������       ��G�����?�            `i@r      s                   �?�6����?a            @b@������������������������       ��LQ�1	�?             7@������������������������       �ד�w��?Q            �^@u      x                   �?�G��l��?            �x@v      w                   �?���1�?s            �f@������������������������       �                      @������������������������       ��.�8�?n            �e@y      z                   �?r�����?�            @k@������������������������       ����7�?             F@������������������������       ��;Eq���?p            �e@|      �                   �?��˶��?�           ��@}      �                   �?������?7            �T@~      �                    �?������?             ;@      �                   �?ףp=
�?             $@������������������������       �r�q��?             @������������������������       �                     @�      �                   �?ҳ�wY;�?
             1@������������������������       �                     "@������������������������       �      �?              @�      �                    �? �Jj�G�?&            �K@�      �                   �?���7�?             6@������������������������       �                     @������������������������       ��}�+r��?             3@������������������������       �                    �@@�      �                    �?��%}*��?�           h�@�      �                   �?N-Xy�2�?�             v@�      �                   �?8S��U\�?�            `n@������������������������       �gO�~k�?b            @d@������������������������       �X�<ݚ�?0            @T@�      �                   �?��_����?L            �[@������������������������       �¦	^_�?             ?@������������������������       ����Q��?6             T@�      �                   �?���#�?�            �r@�      �                   �?�E��
��?l            �c@������������������������       ���c:�??             W@������������������������       �     x�?-             P@�      �                   �?��g�ao�?Z            �a@������������������������       �~|z����?!            �J@������������������������       �Hg����?9            �V@�      �                   �?�|����?           �@�      �                   �?�g�t+�??           "�@�      �                   �?�=��>u�?�           ��@�      �                   �?���?�           (�@�      �                   �? 5x ��?           �z@�      �                    �?8���!��?�            Pt@������������������������       � ��֛�?\            @b@������������������������       �К�m(ܵ?n            `f@�      �                    �?@�n���?:            �Y@������������������������       �@3����?             K@������������������������       �                    �H@�      �                    �?&<�ރ��?�            �u@�      �                   �?�q�qT�?             h@������������������������       �������?J            @Z@������������������������       �>���Rp�?5            �U@�      �                   �?$M����?\             c@������������������������       �j�*�'�??            �Y@������������������������       � �o_��?             I@�      �                   �?�|(:��?�            �r@�      �                    �?H�!b	�?i            @d@������������������������       ���+��<�?:            �U@������������������������       �`-�I�w�?/             S@�      �                    �?|��Q��?O            �`@������������������������       �     ��?*             P@������������������������       �����X�?%            �Q@�      �                    �?Ч퟈��?�           ��@�      �                   �?�q��:�??           �@������������������������       ���}� �?"           }@�      �                   �?�.6��-�?            }@������������������������       �t��%�?�            �l@������������������������       �ȵHPS!�?�            @m@�      �                   �?��@`r�?i           �@������������������������       �y�^���?#           0}@�      �                   �?�Ś{0��?F            @������������������������       ��7��d��?�            `m@������������������������       �`��F:u�?�            Pp@�      �                   �?8Y�tp��?�          �>�@�      �                   �? �f+j}?&           �@�      �                    �?��c��?�           ��@�      �                   �? 
����w?�           H�@������������������������       ���B��{?d           x�@������������������������       �        9            �V@�      �                   �? UQ\R��?           X�@������������������������       � M��~?�            �@������������������������       ��}��L�?Y            �b@�      �                    �? {L(w?�           �@������������������������       � �<��>�?           �{@������������������������       ����1��p?r            �@�      �                   �?p���r�?�           {�@�      �                   �?���"e�?/           �@�      �                    �?"/<#!�?           �{@������������������������       �>���K[�?p            �g@������������������������       ��;����?�            p@�      �                   �?Z��L��?           Pz@�      �                    �?�+Fi��?B             W@������������������������       ��G�z��?             D@������������������������       �����3��?$             J@�      �                    �?p��2;�?�            �t@������������������������       �\�����?U            �`@������������������������       �D��f*��?            �h@�      �                   �?XG�b��?�           �@�      �                   �?��<D�m�?y           �@�      �                    �?���}��?           ,�@������������������������       �ȑ�zA��?           p�@������������������������       ���7)^Ȼ?�           t�@�      �                    �?���=)�?n           H�@������������������������       �X�s����?�            �j@������������������������       ��Y�ɖ�?�            Pu@�      �                    �?P�i0(�?           H�@������������������������       ���ݾ���?�           �@������������������������       �`�����?:           �@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B�      ���@    ���@     3�@     ,�@    ��@     �@     �@     �@      �@     @     �@     @     ��@      @      }@     �~@      x@     �t@     �k@     �l@     �d@      Z@      T@     �c@     �_@      @     �X@              <@      @      3@      �?      3@                      �?      �?             �g@      *@     �g@      "@     �a@       @     �W@       @      W@       @      W@                       @       @             �G@             �G@      @     �G@                      @      @      @      @                      @     ��@     �@     ��@     x�@     l�@      b@     P�@     �Z@     0�@     �G@       @              �@     �G@     ��@     �G@     �@     �B@     p�@      =@     0s@       @      >@      $@     @Q@             �v@     �M@      u@      M@      @             �t@      M@     ps@      D@      j@      @@     �Y@       @      6@      2@      >@      �?      (@      �?      2@              @     �C@              9@      @      ,@      @      @      @      @      @      @      �?      @      �?      @              @    �B�@     ��@     f�@     0~@     ��@      r@     F�@      V@     �@      @     �@      @     В@             ��@     �T@     @�@     �G@     ��@      B@      w@      i@     �l@     @Z@     @a@     �W@     `�@     `h@     �@     �U@     ��@      @     8�@      @     �@             ��@      T@     ��@      ?@     ��@     �H@     pr@     @[@     �f@     �G@     �\@      O@     ��@     �M@     (�@      :@     {@      ,@     @g@      @     �n@      &@     @q@      (@     @V@             `g@      (@     �V@     �@@     �J@      .@     �B@      2@     @w@     h�@      k@     ��@     �e@     ��@     �Z@     h�@     �O@     �l@      *@      ]@      I@     �\@      F@     pv@     @P@     Pv@     �C@     �]@              J@     �C@     �P@      :@     �m@      F@      f@      3@      E@      @      3@      .@      7@      9@     �`@     �c@     ��@     �`@     @�@     �S@     �{@      @     @Z@     �R@     Pu@      D@     �S@      A@     `p@     �L@     @m@      A@      P@      @     �D@      >@      7@      7@     @e@      5@      j@       @     �H@      3@     �c@       @      <@      &@     ``@     ^�@     J�@     ��@     `�@      �@     x@      0@     @`@      0@     @X@      $@     @X@      "@     �W@      @      2@      @     @S@      �?       @      �?      �?              �?      @                     �@@     ��@     �o@     �|@     �V@     �x@      P@      S@      N@     �H@     �J@      ;@      @      t@      @     �i@      @      ]@             �O@      ;@      "@      ;@      K@             �v@     �d@      R@     `c@     �O@     @Z@     �I@     �U@      (@      3@      "@      I@     r@      "@     `o@      @      f@      @     �R@       @      C@      @     L�@     �t@     ��@     �e@      .@      =@      &@      *@      &@                      *@      @      0@      @              �?      0@     �@      b@     ��@      J@      @             ��@      J@     w@      8@     x@      <@     �i@     @W@     �X@      F@      [@     �H@     �@     �c@     @�@     �J@      :@      �?       @              2@      �?       @      �?      $@             p�@      J@     �x@      >@     �j@      5@     �f@      "@     Pv@      6@     �e@      "@     �f@      *@      g@      Z@      X@     �D@      M@      2@              @      M@      ,@      C@      7@               @      C@      .@     @V@     �O@      E@      ;@              @      E@      5@     �G@      B@              (@     �G@      8@     �u@     ��@      (@     ��@             @b@      (@     �@       @     �|@      �?     �f@      �?     Pq@      $@     �w@      @     �c@      @     �E@      @     �\@      @     `k@      �?     �J@       @     �d@     �t@     
�@     `m@     H�@     @a@     �n@      J@     �[@      A@     �S@      2@      @@     �U@      a@      O@     �Z@      8@      >@     @X@     p�@     �L@     ��@      B@     �u@               @      B@     �u@      5@     py@              @      5@      y@      D@     pr@      6@     �b@      2@     `b@              @      2@      b@     @X@     ��@              .@     @X@      �@     �N@     �Z@      <@     �H@     �@@      M@      B@     ȃ@      .@      n@      5@     �x@     ̹@     ��@     ��@     ��@     k�@     �@     ��@     ��@     ��@     Њ@     ��@     �a@      �?      @     ܓ@      a@     x�@     �X@     @e@     @U@     �\@     �C@      L@      G@     (�@      *@     �t@       @     �q@      @     �~@     �C@     ps@      7@      H@      6@     pp@      �?      f@      0@      2@      0@     �c@             �z@     p�@     �m@      i@      d@     �f@      =@     @f@     �`@       @     @S@      5@      $@      3@     �P@       @     �g@     (�@     �a@     �}@      5@     �}@     @^@      @      H@     �C@      $@     �B@      C@       @     �p@      y@      A@     �x@      1@     �J@      &@      3@      @      A@      1@     pu@      @     @T@      &@     `p@     �l@      @      ^@       @     �S@       @      E@             �[@       @     �I@       @      N@             |�@     �q@     ��@     �b@     ��@      V@      &@       @      @       @      @             `�@     �U@     ��@     @P@     �z@     �D@     `z@      8@      c@      5@     @�@      O@      .@      @      &@      @      @      @      @      �?      @             ȅ@      M@      v@      A@     �u@      8@      o@      0@      X@       @     ��@     �`@     8�@      I@      2@      @      ,@      @      "@       @      @      �?      @             ��@     �G@     q@      ?@     @r@      0@     @]@      @     �e@      "@     ��@     �T@      =@      "@      .@       @      (@      @      @      @      ,@      �?     ؄@     �R@     �q@      G@     �w@      <@     �b@      (@      m@      0@     ��@     �@     Px@     @w@     �f@     �f@      \@      Z@       @      &@     �[@     @W@      Q@     �S@      @      4@     @P@      M@      j@     �g@      \@     @Q@               @      \@     �N@     @X@     @^@       @      E@     �W@     �S@     y@     �t@       @     �R@      @      4@      �?      "@      �?      @              @      @      &@              "@      @       @      �?      K@      �?      5@              @      �?      2@             �@@     �x@     @p@     `k@     �`@     �b@     �W@      Z@      M@     �F@      B@     �Q@     �D@      6@      "@      H@      @@     �e@     @_@     @W@     �O@      K@      C@     �C@      9@     @T@      O@      <@      9@     �J@     �B@     X�@    �a�@     �r@     Ф@     @d@     X�@     @Y@      �@      (@      z@      &@     �s@      @     �a@       @     `e@      �?     �Y@      �?     �J@             �H@     @V@      p@     �H@     �a@      <@     @S@      5@     �P@      D@     @\@      :@     @S@      ,@      B@     �N@     `m@       @     @c@      @     �T@      @     �Q@     �J@     @T@     �@@      ?@      4@      I@     �`@     t�@      S@     ��@      ;@     `{@     �H@     �y@      6@      j@      ;@     �i@     �M@     @�@      8@     �{@     �A@     �|@      7@     �j@      (@      o@     �@    �-�@      (@     �@       @     ܝ@       @     8�@       @     h�@             �V@      @     @�@      @     �@       @     �b@      @     ��@       @     �{@       @     �@     ��@     e�@      r@     �@      a@     `s@      D@     �b@      X@      d@      c@     �p@     �B@     �K@      2@      6@      3@     �@@     �\@     �j@     �H@     �T@     �P@     ``@     �n@     "�@     �c@     ��@      ^@     L�@      J@     Ї@      Q@     d�@      B@     (�@      .@     �h@      5@      t@     �V@     (�@      9@     H�@     @P@     �@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r   h%�r  Rr  (KM��r  hm�BXh         J                   �?��0o���?�e           �@       �                    �?F��� \�?#M           l�@       �                    �?� z
��?�3          �Y�@       E                    �?��R%��?�$           ��@       4                    �?���RKN�?�           �@                           �?�dU%�r�?�           �@                           �?ȅ�.��?k           �@                            �?�ȉ5��?f           ��@	       
                     �?V�r��?�           ؇@������������������������       ����f��?           0~@������������������������       �d.��i�?�            �q@������������������������       �:\��M7�?�            �o@                           �?"pc�
�?             &@������������������������       �                     @������������������������       �      �?             @       %                    �?X[+��&�?�           �@                           �?�������?_           _�@                           �?���[�ڥ?�            0q@                            �? =[y��?V             a@������������������������       �����q�?C            @[@������������������������       �PN��T'�?             ;@������������������������       �        T            `a@                           �?�w� `l�?�           L�@                            �?x�}b~|�?+           ��@                           �?8����?�           ��@������������������������       �P�ؑ>�?s           ��@������������������������       ��q�q�?             8@                           �?��L~1_�?�            0p@������������������������       ��R�� �?�             n@������������������������       ��X�<ݺ?             2@       "                    �?aB����?�	           �@        !                     �?��< ���?�           $�@������������������������       ��Qv���x?Y           ��@������������������������       ����m7�?�           (�@#       $                     �?���	�޹?�           ��@������������������������       � ʋ�7�?�           Б@������������������������       �ػn�|Ź?�           ��@&       -                     �?�Z��?4           ̚@'       *                    �?�ʈD��?e           �@(       )                    �?8���lR�?1           p~@������������������������       ������?X            �b@������������������������       ����͡?�            0u@+       ,                    �?ܚI���?4           `@������������������������       �      �?              @������������������������       ��c�L��?.           �~@.       1                    �?dU�oT�?�           ��@/       0                    �?��
Bo5�?�            �v@������������������������       ��q�q��?:             X@������������������������       ���,6"Ѣ?�            �p@2       3                    �?�CV��?�            �v@������������������������       ������H�?             "@������������������������       �������?�             v@5       >                    �?F;w����?�           ��@6       7                    �?jQ��?@           P�@������������������������       �                     $@8       ;                    �?    �\�?;            �@9       :                     �?��(\���?�             n@������������������������       ��8��8��?Y             b@������������������������       �      �?=             X@<       =                     �?|�l�]V�?�             q@������������������������       �Fmq��?b            �c@������������������������       ��d�
t��?C            @\@?       B                    �?,�59�|�?L           �@@       A                     �?�8��Vɯ?�            pu@������������������������       ��g<a�?Z            @c@������������������������       � 7���B�?s            �g@C       D                     �?<5�����?            �h@������������������������       ��/e�U��?E            �[@������������������������       �JyK���?:            �U@F       c                     �?�j����?           ��@G       X                    �?ܺ����?           ��@H       S                    �? )�j��?�           L�@I       N                    �?@i����?�           ��@J       M                    �?`�21�?�            �u@K       L                    �?      �?N             `@������������������������       �      �?             8@������������������������       �      �??             Z@������������������������       ����\=y�?�             k@O       R                    �?0�����?�            �s@P       Q                    �?���̅ӟ?x            �g@������������������������       �                     @������������������������       ��b��fl�?t             g@������������������������       �PF��t<�?^            �_@T       W                    �? +NU�ce?�           �@U       V                    �?@����?�             j@������������������������       �                     7@������������������������       ��1�:2�?y            @g@������������������������       �        [           `�@Y       ^                    �?�Дc3��?y           �@Z       ]                    �?�[�(�V�?O           �~@[       \                    �?��k��?            x@������������������������       �                     5@������������������������       ����(-�?�            �v@������������������������       ��کd�?H            �Y@_       b                    �?>�ܡN��?*           �}@`       a                    �?,I�e���?�            �r@������������������������       ��8��8��?             (@������������������������       �p�z���?�             r@������������������������       ��&�+�?m            `e@d       y                    �?�Œ��?�           Z�@e       n                    �?X�â�?o            �@f       k                    �?`/!}�p�?�           �@g       j                    �?���+�?�            �k@h       i                    �?^��YY��?�            `j@������������������������       ��ӖF2��?/            �Q@������������������������       �:�.���?U            �a@������������������������       �                     &@l       m                    �?�N[��?.           P~@������������������������       �`F	W��?(           �}@������������������������       ����!pc�?             &@o       t                    �?��ѿ�A�?�           ��@p       s                    �?(;L]n�?�            �t@q       r                    �?`��7�ѝ?|            `i@������������������������       �                      @������������������������       ��\=lf�?{             i@������������������������       ���b�h8�?O            �_@u       x                    �?/4���?�           ��@v       w                    �?��wU��?
           y@������������������������       �                     �?������������������������       ��ڊ�e��?	            y@������������������������       �t?�%�y�?�             v@z                           �?�C��2(�?�           ��@{       ~                    �?Ȝw{e��?[           x�@|       }                    �?���.�*�?�            �u@������������������������       �        3             V@������������������������       �P����u�?�             p@������������������������       ���yG���?t            �f@�       �                    �?�	a�$a�?3           x�@������������������������       � !ַЕw?�           <�@������������������������       �b$Vx��?�            �p@�       �                    �?�[K��?�           ��@�       �                     �?�\'PH�?q           x�@�       �                    �?P����?�            �@�       �                    �?`�V0�E�?d            �@�       �                    �?djB���?�            �t@������������������������       �                     @������������������������       ��ߪ5�?�            0t@�       �                    �?�5g����?�            @k@������������������������       �z�G�z�?             $@������������������������       ��n_Y�K�?�             j@�       �                    �?(Ԑ����?            �@������������������������       �t�F>s}�?           �y@������������������������       ��^n��m�?           �|@�       �                    �?�p*4�9�?�           В@�       �                    �?��E��?^           0�@�       �                    �?�ͧJ{�?�            �l@������������������������       ����Q��?             $@������������������������       ��	3��?�            `k@�       �                    �?$	4�}�?�            t@������������������������       �                     @������������������������       ����C��?�            �s@�       �                    �?�
�y�?�           p�@�       �                    �?`�JBjH�?j            �d@������������������������       �                     &@������������������������       ��n_Y�K�?b            �c@������������������������       ���_��	�?'           p~@�       �                     �?n;�]1�?z           ت@�       �                    �?d9��H��?�           @�@�       �                    �?��-���?V           x�@�       �                    �?+�M��?R            �`@������������������������       �                     *@������������������������       �H�tL��?K            @^@�       �                    �?HP�s��?           �z@������������������������       �                     @������������������������       �č��m�?           0z@�       �                    �?�`TV���?H           �@�       �                    �?�ٍ���?M             ]@������������������������       ��S����?             3@������������������������       ��W*��??            @X@������������������������       ���O��[�?�           h�@�       �                    �?�bm��Q�?�           p�@�       �                    �?)O���?�            �v@�       �                    �? ��WV�?!             J@������������������������       �                     $@������������������������       ����N8�?             E@�       �                    �?*-ڋ�p�?�            @s@������������������������       �@�j���?R            @_@������������������������       �^<wr���?y            �f@�       �                    �?����̺?�           И@������������������������       �                     @�       �                    �?����R�?�           ��@������������������������       �     x�?�             x@������������������������       ��{�w�?�           ��@�                          �? ��R�P�?�           %�@�       �                    �?<��}���?}           ��@�       �                    �?������?           ��@�       �                     �?0ڣ-Lͷ?P           ��@�       �                    �?�k.L'>�?�           ��@������������������������       �        '            �N@�       �                    �?�Y�e?�           ~�@�       �                    �? '��h�?�            pt@�       �                    �?      �?�             t@������������������������       ������s�?�            �q@������������������������       �                    �B@������������������������       �����X�?             @�       �                    �?@xF�?�           �@�       �                    �?�ݹ��u�?           �@������������������������       �        �           �@������������������������       �p�<�R�?<           @�@������������������������       �ҳ�wY;�?�            �m@�       �                    �?��@t;}�?�           �@�       �                    �?��y눲�?A           |�@�       �                    �?,(��?R            �_@������������������������       �                     @�       �                    �?������?O            �^@������������������������       �0G���ջ?C             Z@������������������������       �                     3@�       �                    �?hV����?�           ��@������������������������       �                     3@�       �                    �?���~b�?�           4�@������������������������       ���+{�q?,           �|@������������������������       �hl��f�?�           �@�       �                    �?^K�2��?h            `d@������������������������       �                     @������������������������       ��G�z�?f             d@�       �                    �?,�����?�           ��@�       �                    �?Ɔdq��?W            `a@�       �                    �?��a�n`�?O             _@�       �                     �?��M9�U�?D            �[@������������������������       �<�A+K&�?-             S@������������������������       �^������?            �A@�       �                     �?�θ�?             *@������������������������       �      �?              @������������������������       �z�G�z�?             @�       �                     �?�r����?             .@������������������������       �      �?              @������������������������       �                     @�       �                    �?l-MIڼ�?`           |�@�       �                     �?�&/�E�?�           p�@�       �                    �?,�`@��?�           0�@������������������������       ��g���~?�            �p@������������������������       �Tىq��?           �{@�       �                    �?��d5z�?           `y@������������������������       �@��<W��?d            �c@������������������������       �� � J��?�            �n@�       �                     �?���v��?�            0p@������������������������       �B�F<��?b             c@������������������������       ���J���?C            �Z@�       �                    �?��Д?L�?v           \�@�       �                    �?@Q����?,           |@�       �                    �?�B:�g�?u            �e@�       �                    �?@�z�G�?5             T@������������������������       �                      @�       �                     �?�(�Tw�?3            �S@������������������������       �                    �B@������������������������       ���Y��]�?            �D@������������������������       �        @            �W@�       �                    �?إ���?�            0q@�       �                     �?ڇ����?f            @b@������������������������       ��q�q��?C             X@������������������������       ����Q��?#             I@�       �                     �?�+��0��?Q             `@������������������������       �����?4            @S@������������������������       �      �?             J@�                          �?��ݡ�?J           ��@                           �?�S�z��?           p{@������������������������       �ĭ����?�            @o@������������������������       �8����?x            �g@                          �?��+����?,           �}@������������������������       �|�űN�?�            @m@������������������������       ����0���?�            �n@      3                   �?�(@B��?&           ��@                         �?��7e�x�?           (�@      	                   �?�a$��?!           �@������������������������       �                     @
                         �?�5+3���?           ��@                         �?�GA����?�           �@                          �?�*�w�?�             n@                         �?��S�ۿ?Z            �`@������������������������       ����"͏�?            �B@������������������������       �        B            �X@                         �?�iʫ{�?H            �Z@������������������������       �����"�?             =@������������������������       �        2            @S@                         �?(��6�ռ?            {@������������������������       �                      @                          �?��$xtW�?           �z@������������������������       �T�y���?�            `j@������������������������       �0zAA�ڸ?�            �j@                         �?�4�����?c            `c@������������������������       �                     @                          �?�z�G��?_            �b@������������������������       ���Q���?1             T@������������������������       �L�w�=�?.            �Q@      ,                   �?~[���?^           8�@      %                   �?�q�Q�?            ~@      "                   �?0,Tg��?-             U@       !                    �?�~t��?%            @Q@������������������������       �H%u��?             9@������������������������       �fP*L��?             F@#      $                    �?z�G�z�?             .@������������������������       ��q�q�?             @������������������������       �r�q��?             (@&      )                    �?�8��8��?�            �x@'      (                   �?���ȑ��?�             j@������������������������       �        "             N@������������������������       �l������?^            �b@*      +                   �?h�O,��?n            `g@������������������������       ��#-���?            �A@������������������������       �h�˹�?X             c@-      0                   �?D;����?C            �Y@.      /                    �?�q�q�?             .@������������������������       �                     @������������������������       ��eP*L��?             &@1      2                    �?�eP*L��?<             V@������������������������       �`՟�G��?             ?@������������������������       �F�����?"            �L@4      =                    �?�,�9T�?�           �@5      6                   �?�؜�K=�?�           ��@������������������������       �        X             a@7      :                   �?�G�	F��?>           `�@8      9                   �?3k���?C            @\@������������������������       �����X�?&            �O@������������������������       ����H.�?             I@;      <                   �?�w@]D��?�            �y@������������������������       ���p\�?f            �d@������������������������       �$�q-�?�            �n@>      E                   �?I"9k4�?           `�@?      @                   �?     ��?�             r@������������������������       �                     @A      B                   �?ĜA4k�?�            �q@������������������������       �        (             N@C      D                   �?�Cc}h��?�             l@������������������������       �o����?$             M@������������������������       ����O1��?l            �d@F      I                   �?8�NBK��?V           `�@G      H                   �?��SK�?x            �g@������������������������       �����e��?Q            �`@������������������������       ��ݜ����?'            �M@������������������������       �Фղ(k�?�            �t@K      �                    �? #���9�?�           ��@L      }                   �?�q�l�W�?1
           `�@M      p                   �?������?U           �@N      c                   �?�P�
y�?�           $�@O      Z                   �?�j�ߗu�?q           ��@P      W                   �?���_k��?�            v@Q      T                   �?0%*��?�            �k@R      S                   �?� ��1�?            �D@������������������������       �                     �?������������������������       �z�G�z�?             D@U      V                   �?@���=��?q            `f@������������������������       �                     @������������������������       ��B:�g�?m            �e@X      Y                   �?�������?I            �`@������������������������       ��4F����?            �D@������������������������       ������?4             W@[      `                   �?�)��S��?�            `n@\      ]                   �?��}���?_            @c@������������������������       �                      @^      _                   �?d1<+�C�?[            @b@������������������������       �<���D�?            �@@������������������������       �����?E            @\@a      b                   �?�x�E~�?;            @V@������������������������       �        !            �I@������������������������       ��}�+r��?             C@d      k                   �?�lO�m�?           ��@e      h                   �?����?)           �@f      g                   �?��	l�?�             t@������������������������       �                      @������������������������       ��������?�            �s@i      j                   �?��KL�6�?q            �g@������������������������       �                     @������������������������       ���<b�ƥ?n             g@l      m                   �?$�ȻU��?�            `w@������������������������       �                     @n      o                   �?h*�'=P�?�            �v@������������������������       �0�#�.^�?r            `g@������������������������       ������H�?v            �f@q      x                   �?Fmq��?�            �s@r      u                   �?|�{���?\            �`@s      t                   �?$�q-�?             *@������������������������       ������H�?             "@������������������������       �                     @v      w                   �?����?T            �^@������������������������       ��k�'7��?&            �L@������������������������       ��G\�c�?.            @P@y      z                   �?n60�F2�?t            �f@������������������������       �                    �A@{      |                   �?���+�?^            �b@������������������������       �$gv&��?$            �M@������������������������       �:��?:            @V@~      �                   �? YJ��?�           ��@      �                   �?@�E�x�?�           p�@�      �                   �?`��@�F�?a             c@������������������������       �                     *@�      �                   �?@4և���?\            �a@������������������������       ���r._�?            �D@������������������������       �Pa�	�?C            �X@�      �                   �? ۔�.��?J           ��@������������������������       �        0            �S@������������������������       � ���ؑ?           p|@�      �                   �?� �PJ��?1           ��@�      �                   �?    �S�??            �@�      �                   �?x疑��?r            `f@������������������������       ��q�q�?             ;@������������������������       ��˹�m��?_             c@�      �                   �?������?�            �t@������������������������       �~X�<��?-             R@�      �                   �?��d�0-�?�            Pp@������������������������       �                      @������������������������       �0_�n~f�?�            0p@�      �                   �?(��Le�?�           ��@�      �                   �?o����?w            �e@������������������������       ����H.�?$             I@������������������������       ��BE����?S             _@�      �                   �?��'>�{�?{           �@������������������������       ���'���?�            �m@������������������������       ��aR�?�           p�@�      �                   �?      �?[           ض@�      �                   �?��.���?�           *�@�      �                   �?}*��@�?�           T�@�      �                   �?�ș�j�?           P|@�      �                   �?X�*2���?           �z@�      �                   �?8�A�0��?*            �P@�      �                   �?f���M�?             ?@������������������������       �                     �?������������������������       ��q�q�?             >@������������������������       �z�G�z�?            �A@�      �                   �?�4$�?�            �v@�      �                   �?h�����?:             U@������������������������       �`2U0*��?             9@������������������������       ����#�İ?*            �M@������������������������       �  
�R�?�            �q@������������������������       �                     6@�      �                   �?ة��'n�?�           @�@�      �                   �? /8��?�            �p@�      �                   �? ���v�?_             a@������������������������       �        A             W@������������������������       �`Ӹ����?            �F@�      �                   �?�U���?N            �_@������������������������       �        '             L@������������������������       �0z�(>��?'            �Q@�      �                   �?�rӴ��?�           @�@�      �                   �?P`���?�            �y@������������������������       ���I�~R�?v            �h@������������������������       ��>����?~             k@�      �                   �?�R����?�            �v@������������������������       ���S�ۿ?D            @Z@������������������������       �@�p��?�             p@�      �                   �?@���?B            �@�      �                   �?��;���q?^           ��@�      �                   �?����q�?E            @[@������������������������       �                     I@������������������������       ����#�İ?(            �M@�      �                   �? �L�#�Y?           �@������������������������       �        �            �k@������������������������       � ���_?�           |�@�      �                   �?�Cƨ%p�?�            �u@�      �                   �?�P�*�?Q             _@������������������������       �����X�?            �A@������������������������       �N֩	%��?;            @V@�      �                   �?bOvj6��?�            �k@������������������������       �`�Q��?             I@������������������������       �Ї?��f�?u            @e@�      �                   �?tG�o7�?p           ��@�      �                   �?�c:��?�             w@�      �                   �?X���[�?`            �b@������������������������       �                     2@�      �                   �?:ɨ��?U            �`@������������������������       ��+$�jP�?#             K@������������������������       ��n_Y�K�?2            �S@�      �                   �?����d�?�            @k@������������������������       �                    �I@�      �                   �?���dv~�?p            �d@������������������������       �:W��S��?1             S@������������������������       �\Ќ=��??            �V@�      �                   �?��%��?�           ��@�      �                   �?�7��?j           H�@�      �                   �?=0�_�?Y             c@������������������������       �                     �?������������������������       ��}�+r��?X             c@�      �                   �?�Wv���?            {@������������������������       �                     @������������������������       ��-�0�?           �z@�      �                   �?h(M�?           (�@������������������������       ��}�+r��?�             s@������������������������       �@����?Z           h�@r  tr  bh�h"h#K �r  h%�r  Rr  (KM�KK�r	  hQ�B�       _�@     ��@    �\�@    ��@    ���@    ���@     Z�@     
�@     w�@     �@     ��@     ��@     ��@     p~@     ��@     P~@      |@     �s@     �o@     �l@      h@     �U@     �T@     @e@      "@       @      @               @       @     ��@     pw@     ��@     �g@     �p@      @     @`@      @     �Z@       @      7@      @     `a@             ��@      g@     `�@     �R@     ��@      B@     �@      ?@      3@      @     �k@     �C@     `i@      C@      1@      �?     �@     �[@     ��@      (@     ��@      @     �@       @     (�@     �X@     ܐ@     �N@     ��@     �B@     �@      g@     �@      W@     �{@     �G@     �Z@     �D@     �t@      @     �|@     �F@      @      �?      |@      F@     Ѓ@      W@     Ps@      K@     �G@     �H@     `p@      @     Pt@      C@       @      �?     �s@     �B@      h@     8�@     �^@     �x@              $@     �^@     Px@      2@     �k@      (@     �`@      @     �V@     @Z@     �d@     �O@      X@      E@     �Q@     @Q@     �}@      &@     �t@      @     �b@      @     �f@      M@     �a@     �A@      S@      7@      P@     z�@     ��@     t�@     ��@     �x@     (�@     �x@     �p@     �T@     pp@      P@      P@      (@      (@      J@      J@      2@     �h@     `s@      @     `g@      @      @             �f@      @     �^@      @      �?     ��@      �?      j@              7@      �?      g@             `�@     ��@     �m@     �y@     �S@     0w@      .@      5@             �u@      .@     �C@      P@     �s@     �c@     �p@      A@      &@      �?     p@     �@@      G@     @_@     ��@     ��@     �@     8�@     �V@     H�@     �O@     �c@      J@     �c@      @     �P@     �G@     @W@      &@              ;@     �|@      3@     p|@       @      @     ��@     �W@     �s@      &@      i@      @       @             �h@      @     �]@       @      �@     �T@     �v@      B@      �?             �v@      B@     0s@     �G@     �d@     �@     @S@      |@      @     Pu@              V@      @     �o@      R@     @[@     �V@     �@      @     0�@     �U@      g@     ��@     ò@     `�@     @�@     pz@     �@      v@     @h@      l@     �Z@              @      l@     �X@     @`@      V@       @       @      `@      T@     @Q@     ��@      D@     0w@      =@     �z@     Pt@     x�@     �i@     �u@     @e@     �M@      @      @     �d@     �K@      B@     �q@              @      B@     �q@     �]@     ��@      X@     �Q@              &@      X@      N@      7@      }@     �@     �@     `l@     ��@     �Z@     @|@     @R@     �N@              *@     @R@      H@      A@     px@              @      A@     x@      ^@     H�@     �J@     �O@      @      0@      I@     �G@     �P@     P�@     `q@     �@     �g@     @e@       @      I@              $@       @      D@     �g@      ^@     �W@      ?@     �W@     @V@      V@     p�@              @      V@     \�@      5@     �v@     �P@     ��@     ڻ@     �@     ��@     l�@     ��@     {@     �@     �k@     �@      ^@     �N@             ��@      ^@     �s@      .@     `s@      $@     q@      $@     �B@               @      @     �@     @Z@     �@      5@     �@             �@      5@     @c@      U@     p�@     �Y@     ��@     �G@     @^@      @      @             @]@      @     �X@      @      3@             ܑ@     �D@      3@             ��@     �D@     �|@      �?     Ȅ@      D@      [@     �K@              @      [@      J@     \�@     `j@     �X@     �D@      X@      <@     �U@      9@     �O@      *@      7@      (@      $@      @      @       @      @      �?       @      *@       @      @              @     Ԓ@     @e@     t�@     �O@     ��@     �C@     �p@      �?     py@      C@     �w@      8@     �c@      �?      l@      7@      c@     �Z@     �S@     @R@     @R@      A@     �e@     ��@     �V@     pv@      �?     �e@      �?     �S@               @      �?     @S@             �B@      �?      D@             �W@     @V@     @g@     �I@     �W@      ?@     @P@      4@      >@      C@     �V@      9@      J@      *@     �C@     �T@     �@     �E@     �x@      :@      l@      1@     �e@      D@     p{@      0@     @k@      8@     �k@     ؔ@     T�@     H�@      o@     ��@     �Y@      @             ��@     �Y@     p�@     �J@     �j@      ;@     �_@      "@      <@      "@     �X@              V@      2@      &@      2@     @S@             �y@      :@       @              y@      :@     �h@      .@     �i@      &@     @Z@      I@              @     @Z@     �F@      M@      6@     �G@      7@     `{@      b@     x@     �W@      6@      O@      $@     �M@      @      6@      @     �B@      (@      @       @      �?      $@       @     �v@     �@@     �h@      (@      N@              a@      (@     �d@      5@      @@      @     �`@      2@     �J@      I@      @      $@              @      @      @      H@      D@      1@      ,@      ?@      :@     �d@     t�@     �Q@     x�@              a@     �Q@     `|@     �C@     �R@      2@     �F@      5@      =@      ?@     �w@      (@      c@      3@     �l@     �W@     p�@     �F@     `n@              @     �F@     �m@              N@     �F@     `f@      5@     �B@      8@     �a@     �H@     �}@     �@@     �c@       @     @`@      ?@      <@      0@     �s@     �@     /�@     L�@     �@     x�@     �v@     x�@     `m@     `z@     �e@     �s@      C@     `j@      "@     �@@       @              �?     �@@      @     @f@      �?      @             �e@      �?      Z@      =@      *@      <@     �V@      �?     �Z@      a@      4@     �`@               @      4@     �_@      @      =@      0@     @X@     �U@       @     �I@              B@       @     ��@     �N@     �~@      6@      s@      2@       @             �r@      2@      g@      @      @             �f@      @     �t@     �C@      @             �t@     �C@      e@      3@      d@      4@      h@     �_@     �U@     �H@      �?      (@      �?       @              @     @U@     �B@     �G@      $@      C@      ;@     �Z@     @S@             �A@     �Z@      E@     �G@      (@     �M@      >@     �f@     H�@      ,@      �@      $@     �a@              *@      $@     @`@      @      A@      @      X@      @     ��@             �S@      @     0|@     �d@     �@     �L@     p|@      5@     �c@      "@      2@      (@     �a@      B@     �r@      3@     �J@      1@     �n@               @      1@     @n@     �[@     ��@     �O@     �[@      5@      =@      E@     �T@     �G@     p�@      .@      l@      @@     p�@     ؖ@     "�@     L�@     �@     (�@     �|@      N@     �x@      C@     �x@      ;@     �C@      4@      &@              �?      4@      $@      @      <@      &@      v@      @     @T@      �?      8@       @     �L@       @     q@      6@             p�@     �P@     0p@      @     �`@       @      W@             �E@       @      _@      @      L@              Q@      @     X�@     �N@     @x@      9@     �g@      "@      i@      0@     pt@      B@     �X@      @     �l@      =@      a@     ܘ@      @     ��@       @     �Z@              I@       @     �L@      �?     �@             �k@      �?     x�@     �`@     @j@      J@      R@      $@      9@      E@     �G@     �T@     @a@      0@      A@     �P@      Z@     0r@     @�@     @g@     �f@      W@      M@              2@      W@      D@      F@      $@      H@      >@     �W@      _@             �I@     �W@     @R@     �C@     �B@     �K@      B@     @Z@     Ԡ@      >@     X�@       @      b@              �?       @      b@      6@     �y@              @      6@     Py@     �R@     ��@      0@      r@     �M@     |�@r
  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h7Kh8Kh9h"h#K �r  h%�r  Rr  (KK�r  hQ�C              �?r  tr  bhEhUh@C       r  �r  Rr  hYKhZh[Kh"h#K �r  h%�r  Rr  (KK�r  h@�C       r  tr  bK�r  Rr  }r  (hKheM�hfh"h#K �r   h%�r!  Rr"  (KM��r#  hm�B�k         H                   �?�#���?xe           �@       �                    �?L2��?�9          ���@                            �?D��xǣ�?b(          ���@������������������������       � �(y��?           �|@       �                    �?X�SJK�?C'          ���@       G                     �?�O�h�
�?r"          ��@       
                    �?h�G�cG�?\          ���@       	                    �?jIp����?�            �p@������������������������       �p�ݯ��?�            �p@������������������������       �                     @       ,                    �?�/�瓴�?�           �@       !                    �? %�7#-�?�           |�@                           �? k͛��?�	           �@                           �?��K2��?�            �q@                           �? ��F�}?�            0q@                           �?�ۘ�E-�?            @i@������������������������       ��q�q�?>             X@������������������������       �        A            �Z@������������������������       �        ,            @R@                           �?����X�?             @������������������������       �                      @������������������������       �                     @                           �? �XWP��?�           ��@                           �?�63�q�?&           P�@                           �?Hn�.P��?           0�@������������������������       ������ݻ?a           P�@������������������������       �������?�            �o@������������������������       �tk~X��?             B@                            �? ��j�'x?�           "�@                           �? �,a�:s?i           �@������������������������       � -�k$��?v           ��@������������������������       �        �           8�@������������������������       ����N��?f            `c@"       '                    �?,mG����?P           8�@#       &                    �?|�U&k�?�            �k@$       %                    �?��3N�?�            �g@������������������������       �������?V             ^@������������������������       ����L��?.            �Q@������������������������       �      �?             @@(       )                    �?�$9�Ɨ?�           H�@������������������������       �@ѽ�֞?�            pt@*       +                    �? �w5�?�             v@������������������������       ����pA�?�            `q@������������������������       ��"w����?1             S@-       <                    �?ر�#��?�	            �@.       3                    �?�dNC��?�           *�@/       0                    �?�|���?�           ��@������������������������       ��C��2(�?             6@1       2                    �?��W�ƹ?�           8�@������������������������       �                     �?������������������������       ��}��F̹?�           4�@4       9                    �?�����?           ę@5       6                    �? �p8#ګ?]           8�@������������������������       �                     @7       8                    �?��#��?Y           (�@������������������������       �                    �B@������������������������       �P������?B           ��@:       ;                    �?��8�$>�?�            0r@������������������������       �                      @������������������������       ��#*�'ʴ?�            �q@=       B                    �?4^�0/�?�           �@>       ?                    �?z�G�z�?             4@������������������������       ��z�G��?             $@@       A                    �?ףp=
�?             $@������������������������       �      �?              @������������������������       �                      @C       F                    �?p�(���?�           ��@D       E                    �?l�6�?C           p�@������������������������       �\�m�Y�?"           }@������������������������       �x��-�?!           �}@������������������������       ��L���?p             g@H       S                    �?���Uf��?           "�@I       J                    �?�nf1���?�            `t@������������������������       ��ՙ/�?�            �l@K       P                    �?�¦�{��?6            �W@L       O                    �?X��Oԣ�?$             O@M       N                    �?     ��?             @@������������������������       ��������?             >@������������������������       �                      @������������������������       �                     >@Q       R                    �?�FVQ&�?            �@@������������������������       �����X�?             @������������������������       �                     :@T       o                    �?��b�h8�?O           ܱ@U       b                    �?.��uo��?k           ��@V       _                    �?�禺f��?�            �x@W       X                    �?��5Վ3�?�            Pv@������������������������       �                     �?Y       \                    �?��Έ�D�?�            @v@Z       [                    �?؇���X�?�            �m@������������������������       �����?�            @l@������������������������       �r�q��?	             (@]       ^                    �?|�9ǣ�?J            �]@������������������������       �����&��?B            �Z@������������������������       �                     (@`       a                    �?�	j*D�?            �C@������������������������       �      �?             @@������������������������       �                     @c       d                    �?�^����?q            �d@������������������������       �                      @e       j                    �?ؓ��M{�?p            �d@f       i                    �?F��ӭ��?d             b@g       h                    �?�s��:��?M            �\@������������������������       �l��[B��?8            �U@������������������������       ��q�q�?             ;@������������������������       �d��0u��?             >@k       n                    �?�����?             5@l       m                    �?      �?             0@������������������������       ��8��8��?             (@������������������������       �      �?             @������������������������       �                     @p                           �?���D�?�	           R�@q       x                    �?P��IV��?�           ܫ@r       u                    �?(2����?�           ��@s       t                    �?���{}�?,           ��@������������������������       ��>���?z           P�@������������������������       � ���v�?�             q@v       w                    �? �-��?�           8�@������������������������       ����N8�?�           ��@������������������������       ����d�?�            �u@y       |                    �?@q���?�           �@z       {                    �?XU�s*P�?�           H�@������������������������       �� ��߈?<           �~@������������������������       ��dD��?�           8�@}       ~                    �?����Ձ�?            {@������������������������       �        _            `d@������������������������       �0M����?�            �p@�       �                    �?@�+�V�?           �{@�       �                    �?�e���@�?d            @c@������������������������       �@uvI��?A            �X@������������������������       ��h����?#             L@�       �                    �? ��s`�?�            r@������������������������       �Pq�����?o            @e@������������������������       �0x�!���?L            �]@�       �                    �?8p9(���?�           Ȟ@�       �                    �?$	4�}�?B            �Z@�       �                     �?�o��gn�?0            �T@�       �                    �?$�q-�?             J@�       �                    �?�?�|�?            �B@������������������������       ��nkK�?             7@������������������������       �                     ,@�       �                    �?z�G�z�?
             .@������������������������       �r�q��?             @������������������������       ��<ݚ�?             "@�       �                    �?��a�n`�?             ?@�       �                    �?�GN�z�?             6@������������������������       ��q�q�?             .@������������������������       �                     @�       �                    �?�<ݚ�?             "@������������������������       ��q�q�?             @������������������������       �                     @�       �                    �? �q�q�?             8@�       �                     �?      �?              @������������������������       �r�q��?             @������������������������       �                      @������������������������       �                     0@�       �                     �?��B��?�           �@�       �                    �?r��Xo�?�           8�@�       �                    �?��d�H2�?�           h�@�       �                    �?�q5���?{           ��@������������������������       ������?�            �v@������������������������       ��~����?�            �m@������������������������       �r�q��?#             K@�       �                    �?�7a��r�?           |@�       �                    �?6]�f!��?�            0v@������������������������       ���E���?v            �h@������������������������       ��;u�,a�?d            �c@������������������������       �,�[I'��?8            �W@�       �                    �?pu+xi �?�           ȇ@�       �                    �?�/�L���?�            @w@������������������������       ��W;�E��?�            �j@������������������������       �v�_���?^            �c@�       �                    �?=q�$��?�            Px@�       �                    �?��@C'�?�            `l@������������������������       �x����6�?d             c@������������������������       �������?-            �R@�       �                    �?      �?h            @d@������������������������       �X�����?<             V@������������������������       ���+��?,            �R@�       �                     �?4�	~���?�           û@�       �                    �?x^:��K�?�           ��@�       �                    �?��c:�?�           @�@�       �                    �?x*pY1��?\           h�@�       �                    �?�Ws�x��?�            �i@�       �                    �?�c�Α�?             =@������������������������       ����|���?             6@������������������������       �                     @�       �                    �?t�#�$�?p             f@�       �                    �?��^@=��?Y            ``@������������������������       �ܐ҆��?>            @W@������������������������       �P����?             C@������������������������       ����.�6�?             G@�       �                    �?|�űN�?�            �u@�       �                    �?85�}C�?�            �n@������������������������       �X�s����?�            �j@������������������������       �     ��?             @@������������������������       �PԱ�l�?<            �Z@�       �                    �?�`ص���?_           �@�       �                    �? ��OC�x?�            �t@�       �                    �?��S����?q            �g@������������������������       �                     @������������������������       ���W��#�?l             g@������������������������       �        c            `a@�       �                    �?�HGݐ\�?�            `k@������������������������       �XB���?M             ]@������������������������       �        >            �Y@�       �                    �? �gb��?�           �@�       �                    �?@d���?j           ��@�       �                    �?Pa�.l�?(            �P@�       �                    �?�8��8��?             8@������������������������       �                     3@������������������������       ����Q��?             @�       �                    �?�T|n�q�?            �E@������������������������       �$�q-�?
             *@������������������������       �z�G�z�?             >@�       �                    �?Rt_鏖�?B           ��@�       �                    �?0�I��8�?6            @������������������������       �7��?�            �w@������������������������       �@��,*�?E            �]@�       �                    �? �x���?           0z@������������������������       �D��*�4�?�            @q@������������������������       �d��G,�?W            �a@�       �                    �?4�e��&�?�           ܐ@�       �                    �?��~R���?&            �O@�       �                    �?HP�s��?             9@�       �                    �?@4և���?             ,@������������������������       �                     @������������������������       �؇���X�?             @�       �                    �?�C��2(�?             &@������������������������       �      �?              @������������������������       �                     @������������������������       �                     C@�       �                    �?��tM��?l           ��@�       �                    �?�{����?8           X�@�       �                    �?X�Հ�+�?�            Py@������������������������       ��&=�w��?�            �p@������������������������       ����2���?[            �a@�       �                    �?P&��?I            �]@������������������������       ��Y�R_�?-            �Q@������������������������       ���C���?            �G@�       �                    �?����0�?4           �~@�       �                    �?�:g�1��?�            pv@������������������������       ����?a            �c@������������������������       ��(��?             i@�       �                    �?pб����?T            �`@������������������������       �Ȩ�I��?            �J@������������������������       �gO�~k�?5            @T@�       %                   �?��}*_��?�	           ̮@�                          �?��Љ��?Z           �@�       	                   �?:ª�d�?�            pv@�       �                    �?4;����?�            �p@�       �                    �? qP��B�?7            �U@������������������������       � Df@��?5            �T@������������������������       �                     @�                          �?*;L]n�?�            �f@                          �?:%�[��?f            �a@                         �?&X�IN�?\             `@������������������������       ��0u��A�?W             ^@������������������������       �                     "@������������������������       �$�q-�?
             *@                         �?D�n�3�?             C@                         �?<=�,S��?            �A@������������������������       ��P�*�?             ?@������������������������       �                     @������������������������       �                     @
                         �?��r
'��?D            @W@                         �?xdQ�m��?:            @T@������������������������       � �Cc}�?             <@������������������������       ��&=�w��?(            �J@                         �?�q�q�?
             (@������������������������       �                     @������������������������       �                     @                          �? ~�����?]           ��@                         �?H�te�?�           `�@                         �?`���z[�?�            pt@                         �?p�C��?�            q@������������������������       �                     �?                         �?�����?�             q@������������������������       �0���ަ?l            �e@������������������������       �`�E���?1            @X@������������������������       ��>����?!             K@                         �?썐�b��?�           ��@������������������������       �                     @                         �?tPx���?�           h�@������������������������       ���|�#��?�            0x@                         �?�实HW�?�            �x@������������������������       ��0p<���?w             h@������������������������       �8?W���?�             i@!      "                   �?�q�q�?�            �p@������������������������       �>�`���?T             a@#      $                   �?b �y��?R            �_@������������������������       ��^���U�?%            �L@������������������������       �">�֕�?-            �Q@&      1                   �?���n��?o           >�@'      ,                   �?Z�����?�           t�@(      )                   �?�nkK�?G           �@������������������������       ������?1           P}@*      +                   �?$G$n��?            �B@������������������������       ��q�q�?             @������������������������       �l��\��?             A@-      0                   �?v��8�?�           �@.      /                   �?�ƶC5{�?-           �~@������������������������       �@A��q�?X            �`@������������������������       �R���Q�?�            �v@������������������������       ��K����?n            �f@2      9                   �?���}���?�           �@3      6                   �?2\Q��?�            Py@4      5                   �?��X
��?�            ps@������������������������       �r֛w���?             ?@������������������������       �P���Q�?�            �q@7      8                   �?`Ql�R�?;            �W@������������������������       ��?�|�?            �B@������������������������       �0�)AU��?#            �L@:      A                   �?|�f���?�           h�@;      >                   �?䯦s#�?#            �J@<      =                   �?8�Z$���?	             *@������������������������       �      �?              @������������������������       �                     @?      @                   �?R���Q�?             D@������������������������       ��z�G��?             $@������������������������       ���S�ۿ?             >@B      E                   �?�ˡ�5��?k           ��@C      D                   �?�Y���?�            �j@������������������������       �\���(�?k             d@������������������������       ���B����?             J@F      G                   �?d��o�t�?�            @v@������������������������       ������?�            �p@������������������������       ��O�w���?:            �V@I      �                    �?�n��o��?�+          �Z�@J      g                   �?���7i��?�           ��@K      X                   �?�����?           ��@L      S                   �?�Pݶ�C�?G           p@M      R                   �?4և����?�             l@N      Q                   �?�IQu`�?u            �f@O      P                   �?$�q-�?_            �a@������������������������       �                     �?������������������������       �,�d�vK�?^            �a@������������������������       �                    �B@������������������������       ��������?             F@T      U                   �? Dl��?�            pq@������������������������       �`�V���?m            �c@V      W                   �?��v$���?O            �^@������������������������       ��Ń��̧?             E@������������������������       �@�z�G�?0             T@Y      d                   �?@c��-�?�           ��@Z      ]                   �?�k~X��?�            �v@[      \                   �?@����?|             j@������������������������       �                     8@������������������������       � S5W�?p             g@^      a                   �?p�`Bh�?e            �b@_      `                   �? ���J��?            �C@������������������������       �                     �?������������������������       �P�Lt�<�?             C@b      c                   �?������?J             \@������������������������       �                     @������������������������       ���?^�k�?G            @Z@e      f                   �? :|�&e\?�           �@������������������������       � �K��l?r           @�@������������������������       �        i           ȁ@h                         �?P��U=�?�           е@i      p                   �?��滵i�?�           |�@j      m                   �?4s��1�?�           ��@k      l                   �? |�'t�?�            @p@������������������������       ������?a             c@������������������������       ��q�q�?G             [@n      o                   �?0��0GY�?(           X�@������������������������       ���~����?�            �x@������������������������       �p��E�m�?5           �}@q      x                   �?P�-8��?�           <�@r      u                   �?f>�cQ�?�           ��@s      t                   �?��	�l��?v            �f@������������������������       �v�X��?=             V@������������������������       �z�J�?9            �W@v      w                   �?|O/(y��?M           0�@������������������������       �|�l�]�?�             q@������������������������       ���ׄ��?�            `q@y      |                   �?��n��?8           0@z      {                   �?�S����?             j@������������������������       ��f7�z�?             =@������������������������       ��?�P�a�?l            �f@}      ~                   �?��1���?�             r@������������������������       ���}*_��?%             K@������������������������       � ,��-�?�            �m@�      �                   �?���Ӧ��?�           $�@�      �                   �?(}t�3_�?r           x�@�      �                   �?�SrN��?�            @o@������������������������       ��e�,��?I            �]@�      �                   �?�N2�,��?N            �`@������������������������       �f�<�>��?#            �M@������������������������       �P�t��?+            @R@�      �                   �?Hv�G�?�            Pu@�      �                   �?X�d1���?�            `l@������������������������       ���|\�d�?l            �e@������������������������       �^(��I�?%            �K@������������������������       ��5C�z�?J            �\@�      �                   �?���DA�?z           ��@�      �                   �?��#��?�           �@�      �                   �?�g+��@�?�           �@�      �                   �?����?�             x@������������������������       �                     �?������������������������       ��C��2(�?�            x@������������������������       �p�$ :u�?
           �@�      �                   �?�x+M���?�            �w@������������������������       �ȵHPS!�?d            �c@������������������������       ����=��?�            @l@�      �                   �?     �?�            �@�      �                   �? "��u�?�            �r@������������������������       �                      @������������������������       �8����?�            �r@������������������������       ��푵V�?�           ��@�      �                   �?��#/���?�           ��@�      �                   �?������?           :�@�      �                   �?`�����?�            �@�      �                   �? �����?            |�@�      �                   �?���2/y�?           �|@�      �                   �?�"P��??            �X@������������������������       �                     @������������������������       ����}<S�?:             W@�      �                   �? ����?�            Pv@������������������������       �        '            �N@������������������������       �PL��V�?�            �r@�      �                   �?`�s���?           \�@������������������������       �H��%�^�?l             d@������������������������       ��F���?�           ؐ@�      �                   �? %��$��?�            r@�      �                   �? �q�q�?=             X@������������������������       �                      @�      �                   �?`�q�0ܴ?;            �W@������������������������       ��L���?            �B@������������������������       �0�)AU��?'            �L@������������������������       �        s             h@�      �                   �?�_/Ap|�?E
           z�@�      �                   �?�Q�*B	�?y           ��@�      �                   �?�A�0�^�?�           ��@�      �                   �?h���
�?            `z@������������������������       ��I{A�?>            �X@�      �                   �?�@�{���?�            0t@������������������������       �                      @������������������������       � ˤ���?�            t@�      �                   �?�5*�?�           Ѓ@������������������������       �\Ќ=��?p            �f@�      �                   �?���=��?           @|@������������������������       �                     @������������������������       ��G���?           �{@�      �                   �?����:��?�           �@�      �                   �?TC4] �?W           ��@������������������������       ��9:�l'�?D            @X@������������������������       ��
���x�?            {@�      �                   �?���s�b�?�           ��@������������������������       ��iޤ��?�            �p@������������������������       � �E����?�           h�@�      �                   �?^@��?�           ��@�      �                   �?>vN#�?�            �j@�      �                   �?�������?J             ]@������������������������       �F�����?'            �L@������������������������       �@�r-��?#            �M@�      �                   �?ڡR����?B            �X@������������������������       ��E��
��?"             J@������������������������       ���c:�?              G@�      �                   �?H�*�ݰ�?@           X�@�      �                   �?��_!�?            z@������������������������       �x�kE�?r            `g@������������������������       ��.^��?�            �l@�      �                   �?����[�?>           H�@�      �                   �?����s�?o            �g@������������������������       �                      @������������������������       �4z�_�\�?n            �g@������������������������       �p�u$v��?�            �v@�      �                   �?�U���?�	            �@�      �                   �?bU�\��?[           ȍ@�      �                   �?xE���?�            �k@�      �                   �?z�G�z�?;            @U@������������������������       � �q�q�?!             H@������������������������       ��Gi����?            �B@������������������������       ��>����?Z            �`@�      �                   �?���[�?�           �@������������������������       �                     @@�      �                   �?�ӕ�?�           �@�      �                   �?Pe6�p�?�            �p@������������������������       �������?p            �f@������������������������       �X�Cc�?:             U@������������������������       ��m,Zez�?           P{@�      �                   �?���t�=�?l           ��@�      �                   �? �o-�?�           l�@������������������������       �P����?$            �M@������������������������       ��n�k���?�           ��@�      �                   �?��IO_��?�           ��@�      �                   �?�<��S��?�            @o@������������������������       �"pc�
�?%            �K@������������������������       ��-� �8�?}            `h@�      �                   �?Х-��ٹ?�           ș@������������������������       �`�g�ɦ�?�            �q@������������������������       �(�Ko��?O           L�@r$  tr%  bh�h"h#K �r&  h%�r'  Rr(  (KM�KK�r)  hQ�B�       U�@     ��@    ���@     �@    �D�@     Ȝ@      l@     �m@     ��@     �@     k�@     (�@     ��@     �z@     `e@     �X@      e@     �X@      @            �`�@     �t@     ��@     �`@     x�@     �L@     pq@      @      q@      �?      i@      �?     �W@      �?     �Z@             @R@              @       @               @      @             J�@      K@     ��@      G@     ��@     �C@     P�@      @@     �n@      @      =@      @     �@       @     �@      @     ��@      @     8�@              c@       @     Љ@     @S@      c@     @Q@     �a@     �H@      V@      @@     �J@      1@      (@      4@     �@       @      t@      @     �u@      @     @q@       @     �R@      �?     ��@     �h@     F�@     �\@     ��@      P@      4@       @     @�@      O@      �?             <�@      O@     ��@      I@     ��@      C@      @             ��@      C@     �B@             ��@      C@     pq@      (@       @             �p@      (@     ��@     �T@      0@      @      @      @      "@      �?      @      �?       @             `�@     �S@     p�@      P@     �z@      A@     �{@      >@     @e@      .@     j�@     �{@     �e@      c@      V@     �a@     �U@      "@     �K@      @      9@      @      7@      @       @              >@              ?@       @      @       @      :@             ��@      r@      {@     ``@     0u@     �L@     �s@     �F@      �?             ps@     �F@     �i@      A@     @h@      @@      $@       @     �Z@      &@     �W@      &@      (@              ;@      (@      4@      (@      @             @W@     �R@               @     @W@      R@     �R@     �Q@     �O@     �I@     �F@      E@      2@      "@      &@      3@      3@       @      ,@       @      &@      �?      @      �?      @             �@     �c@     ��@     �a@     `�@     �T@     x�@      *@     �@      "@     �p@      @     $�@     @Q@     ��@      B@     �s@     �@@     �@     �N@     ��@     �D@     �~@      @     �@      C@     �y@      4@     `d@             `o@      4@     �z@      ,@      c@       @     @X@      �?     �K@      �?     Pq@      (@     @d@       @     �\@      @     H�@      �@      (@     �W@      &@      R@      @      H@      �?      B@      �?      6@              ,@      @      (@      �?      @       @      @      @      8@      @      1@      @      $@              @       @      @       @      �?              @      �?      7@      �?      @      �?      @               @              0@     �@     �@     �@     �x@     P|@      i@     �y@     �g@     �o@     @[@     `c@     �T@     �F@      "@     �o@     `h@     �h@     �c@     �Z@     �V@     �V@      Q@     �L@     �B@     �@     �n@     �p@      Z@     �d@      I@      Z@      K@     �n@     �a@     �d@     �N@     �[@     �D@     �K@      4@     @T@     @T@     �F@     �E@      B@      C@     �@     ��@     n�@     0�@     @�@     �|@     �Z@     0|@     �T@      _@       @      5@       @      ,@              @     �R@     �Y@     �Q@      N@      G@     �G@      9@      *@      @     �E@      8@     pt@      4@      l@      .@     �h@      @      ;@      @     �Y@     ��@      @     pt@      �?     �g@      �?      @             �f@      �?     `a@             �j@      @      \@      @     �Y@             ��@     �u@      �@     @f@      =@      C@      6@       @      3@              @       @      @      B@      �?      (@      @      8@     8�@     �a@     @{@      N@     �u@      <@     �U@      @@     0u@      T@      p@      4@     �T@      N@     X�@     �e@      7@      D@      7@       @      *@      �?      @              @      �?      $@      �?      @      �?      @                      C@     ��@     �`@     �|@      O@      x@      5@     �o@      $@      `@      &@     @S@     �D@     �H@      6@      <@      3@     pz@     �Q@     �t@      ;@     `c@      @      f@      7@     �V@     �E@     �C@      ,@      J@      =@     d�@     Ж@     x�@     �z@     �V@     �p@      T@     @g@       @      U@       @     @T@              @     �S@     �Y@      L@     �U@     �K@     �R@      G@     �R@      "@              �?      (@      6@      0@      6@      *@      2@      *@      @                      @      $@     �T@      @      S@      @      9@       @     �I@      @      @      @                      @     �@     �c@     P�@      Q@     �s@      $@     �p@      @      �?             �p@      @     `e@      @     �W@       @      I@      @     ��@      M@      @             ��@      M@     @v@      ?@     �v@      ;@     �f@      &@      g@      0@      f@      V@     @W@      F@     �T@      F@     �A@      6@      H@      6@     P�@     ,�@     ��@     8�@      6@     @~@      1@     @|@      @      @@       @      �?      @      ?@      �@     ``@     P{@      M@     ``@      @      s@      K@     �Z@     @R@     ��@     @z@     �\@     0r@      6@     r@       @      7@      ,@     �p@      W@       @      B@      �?      L@      �?     �~@      `@      4@     �@@      &@       @      @       @      @              "@      ?@      @      @       @      <@     �}@      X@     �e@      C@     `b@      *@      ;@      9@     �r@      M@      n@      8@     �L@      A@     ��@     ��@     �@     �@      >@     �@      8@     �}@      4@     �i@      &@      e@      &@     �`@              �?      &@     ``@             �B@      "@     �A@      @     0q@       @     `c@       @      ^@      �?     �D@      �?     �S@      @     ��@      @     0v@      �?      j@              8@      �?      g@      @     `b@      �?      C@              �?      �?     �B@      @     @[@              @      @     �Y@      �?      �@      �?     8�@             ȁ@      �@     ,�@     `t@     ��@     �b@     Ў@     @T@     `f@     �F@     �Z@      B@      R@      Q@     8�@     �E@     0v@      9@     @|@      f@     x�@      [@     ��@     �L@     @_@      :@      O@      ?@     �O@     �I@     0@      9@     �n@      :@     �o@     @Q@     �z@     �@@      f@      (@      1@      5@     �c@      B@     �o@      4@      A@      0@     �k@     �u@     h�@     �h@     �x@     �V@     �c@      C@      T@     �J@     �S@      8@     �A@      =@      F@     @Z@     �m@      P@     `d@      I@     �^@      ,@     �D@     �D@     @R@     @c@     R�@     �Z@     d�@     @S@     ��@     �A@     �u@              �?     �A@     �u@      E@     Ȉ@      =@     v@      2@     @a@      &@     �j@      H@     ��@      2@     �q@               @      2@     �q@      >@     ��@      �@     M�@     �@     �@      >@     ��@      :@     �@      ,@     �{@       @     �V@              @       @      U@      @     �u@             �N@      @      r@      (@     ,�@      @     `c@      @     ��@      @     �q@      @      W@               @      @     �V@      @      A@      �?      L@              h@      �@     �@     �v@     ڤ@     `e@     ��@     @S@     �u@     �A@      P@      E@     �q@               @      E@     pq@     �W@     ��@      R@     �[@      6@     �z@              @      6@     �z@      h@     ��@     �J@     �}@      7@     �R@      >@     @y@     �a@     h�@      T@     �g@      N@     x�@      c@     $�@     �R@     `a@     �A@     @T@      :@      ?@      "@      I@      D@      M@      5@      ?@      3@      ;@     @S@     ��@      A@      x@      2@      e@      0@     �j@     �E@     �@      7@      e@               @      7@     �d@      4@     `u@     �o@     �@      U@     (�@      ;@      h@      1@      Q@       @      G@      .@      6@      $@     @_@     �L@      �@              @@     �L@      �@     �A@     �l@      @     �e@      >@      K@      6@     �y@     @e@     :�@       @     L�@      �?      M@      @     d�@     @d@     (�@     �R@      f@      $@     �F@      P@     ``@      V@     h�@      3@     �p@     @Q@     8�@r*  tr+  bubhhubh)�r,  }r-  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h7Kh8Kh9h"h#K �r.  h%�r/  Rr0  (KK�r1  hQ�C              �?r2  tr3  bhEhUh@C       r4  �r5  Rr6  hYKhZh[Kh"h#K �r7  h%�r8  Rr9  (KK�r:  h@�C       r;  tr<  bK�r=  Rr>  }r?  (hKheM�hfh"h#K �r@  h%�rA  RrB  (KM��rC  hm�B(f         �                    �?R���v��?�e           �@       �                    �?��e��?�5          ��@       p                    �?0U�#��?�(           ��@                            �?Hp����?$           W�@������������������������       ��4T���?           �z@                           �?l� ߙ�?�"          ��@                           �?^��S�?/           ؋@                           �?ռ�%�?�           �@	       
                     �?
;&����?I           �@������������������������       �R]�8�?�            `p@������������������������       �vz�M1�?�            �n@                           �?�u�w�u�?`            `d@                            �?<���|��?R            @a@                           �?�X�<ݺ?=             [@������������������������       � ѯ��?<            �Z@������������������������       �                     �?������������������������       �r�q��?             >@                            �?`2U0*��?             9@������������������������       �                     4@������������������������       �z�G�z�?             @������������������������       �        �            �k@       A                    �?�W�3�k�?�            ��@       .                    �?���S�ư?          ���@       %                     �?d�����?e           ��@       "                    �?�Cй��?\            �@                           �?����6�?7           @�@                           �? h����?           H�@                           �?�tVV�?^           ��@������������������������       �                      @������������������������       �����j�?\           ��@������������������������       ����m&�?�            Pq@        !                    �?���N8�?%            �O@������������������������       � �Cc}�?             <@������������������������       �                    �A@#       $                    �?�������?%             N@������������������������       � �o_��?              I@������������������������       �                     $@&       +                    �?4�d����?	            z@'       *                    �?,%*�%�?�            @x@(       )                    �?�d�S��?�            �u@������������������������       �س|G��?�            �m@������������������������       �P�Lt�<�?F            �\@������������������������       ���%��?            �B@,       -                    �?(;L]n�?             >@������������������������       ��X�<ݺ?             2@������������������������       �        
             (@/       6                    �?��V4�Ϊ?�          �0�@0       3                     �? ��T�-?�	           ��@1       2                    �? �$ 3_X?�           ��@������������������������       � ��.lpg?}           Е@������������������������       �        \           ,�@4       5                    �?���!IC�?           \�@������������������������       ��Y��oA�?u           (�@������������������������       �        �           ��@7       :                    �?����>�?�
           �@8       9                     �?������?�           0�@������������������������       �pV�g���?�           (�@������������������������       �Нr����?�           �@;       >                    �?����ꣴ?/           ~�@<       =                     �?`,�I��?
           ��@������������������������       ��_:��"�?R           ��@������������������������       �P����?�           �@?       @                     �?�p�#Rǻ?%           P}@������������������������       ��}�+r��?�            �p@������������������������       ��s��=��?            `i@B       Y                    �?xW����?�           z�@C       L                     �?n��$�?           �}@D       I                    �?���}��?�             s@E       H                    �?p��͇�?�            �q@F       G                    �?�|l=#��?�            �m@������������������������       �tݹ��B�?Y            `c@������������������������       �����!�?0            �T@������������������������       ��I� �?             G@J       K                    �?؇���X�?             5@������������������������       �r�q��?             (@������������������������       ������H�?             "@M       N                    �?������?r            �e@������������������������       �      �?              @O       T                    �?.�qd���?p            `e@P       Q                    �?�O6j���?c            �b@������������������������       �^ۈ��.�?:            �V@R       S                    �?l��[B��?)             M@������������������������       ��ʻ����?             A@������������������������       �      �?             8@U       X                    �?��2(&�?             6@V       W                    �?d}h���?	             ,@������������������������       �z�G�z�?             @������������������������       ��<ݚ�?             "@������������������������       �                      @Z       e                    �?x!�?�           ��@[       ^                    �?�Sa��?�           D�@\       ]                     �?��f�ب?�           �@������������������������       ��?�|�?�             w@������������������������       �p�C��?�            q@_       b                    �? ��7ZH�?Q           p�@`       a                     �? ���l�?�            @x@������������������������       � 4^��?�            �m@������������������������       ����=��?e            �b@c       d                     �?@	tbA@�?T            @a@������������������������       ����E�?4            �U@������������������������       ����J��?             �I@f       i                    �?�`T�
\�?�           <�@g       h                     �?��O`��?            x�@������������������������       �|�:��a�?9           �@������������������������       �H�8i��?�            `w@j       m                     �?(���G2�?{            �@k       l                    �?s;!���?�           ؃@������������������������       ��������?!           0{@������������������������       ��ڊ�e��?u             i@n       o                    �?��|Io��?�            Pv@������������������������       ����Ls�?�            @p@������������������������       ��*v��?@            @X@q       �                    �?���y��?�           ��@r       }                    �?�4B.��?�           x�@s       x                     �?b�h�d.�?            �A@t       u                    �?�����?             5@������������������������       �                     (@v       w                    �?�<ݚ�?             "@������������������������       �      �?             @������������������������       �                     @y       |                    �?����X�?             ,@z       {                    �?�q�q�?
             (@������������������������       ��z�G��?             $@������������������������       �      �?              @������������������������       �                      @~       �                    �?�r����?�           ؏@       �                    �?������?M           ȋ@�       �                     �?��wܒ��?U           �@������������������������       ���d@��?�             t@�       �                    �?���N8�?�            �g@������������������������       �                      @������������������������       �ƿ���c�?�            `g@�       �                     �?�S
�T�?�            �w@������������������������       ��3�w�?�             m@������������������������       ��e����?_             b@�       �                     �?�θ�?M            @`@������������������������       ��A+K&:�?,             S@������������������������       �����|e�?!             K@�       �                    �?Z�8��M�?
            �@�       �                     �?��V�I��?�            �w@�       �                    �?ĹER���?�            `j@������������������������       �                     &@������������������������       �"��u���?�             i@�       �                    �?�t��?k            �d@������������������������       �                     $@������������������������       �d��J_��?e            `c@�       �                     �?������?           �z@�       �                    �?tϺFˁ�?�            @o@�       �                    �?h�g%���?o            �e@������������������������       �      �?             @������������������������       ���ƣ��?k             e@�       �                    �?rOP\6�?4            @S@������������������������       �                     @������������������������       ��J�T�?/            �Q@�       �                    �?��۾%d�?n            �e@������������������������       �        
             3@�       �                    �?��$
���?d            `c@������������������������       �(���@��?9            �W@������������������������       �:2vz�M�?+            �N@�       �                    �?����=*�?�           b�@�       �                    �?���?�           <�@�       �                     �?��n
賳?N           �@�       �                    �?���+�ǲ?>           �}@�       �                    �?`�q�0ܴ?�            �q@�       �                    �?��*��?\            `a@������������������������       �                     �?������������������������       �<���|��?[            @a@������������������������       �@Tn�kq�?c            �a@�       �                    �?�==Q�P�?            �g@�       �                    �?��S�ۿ?(             N@������������������������       �                     @@������������������������       �؇���X�?             <@�       �                    �? ����?W            @`@������������������������       �`�q�0ܴ?!            �G@������������������������       �        6            �T@�       �                    �?0z�(>��?           �z@�       �                    �?����} �?�            �t@������������������������       �                      @�       �                    �?�ɢ����?�            0t@�       �                    �?pXg�Ɛ�?�            �o@������������������������       ��==Q�P�?;            �W@������������������������       �(�5�f��?a            �c@�       �                    �?`����֜?.            �Q@������������������������       �      �?             @@������������������������       �                     C@�       �                    �?<����?A            �W@������������������������       �X�EQ]N�?            �E@������������������������       �0G���ջ?$             J@�       �                    �?�Q�w��?_           h�@�       �                    �?�><˖��?�           ��@�       �                    �?���P7��?.           @�       �                     �?r(�܈�?�            pp@������������������������       ��z�G��?h             d@������������������������       �b*0t��?@            �Y@�       �                     �?.��$�?�            @m@������������������������       �bKv���?O            @a@������������������������       �      �?7             X@�       �                    �?b���L��?�            0r@�       �                     �?�G�z��?l             d@������������������������       ���̅��?C            �W@������������������������       ��G\�c�?)            @P@�       �                     �?��N��?O            ``@������������������������       �z\�3�?/            �S@������������������������       ��	j*D�?              J@�       �                     �?�KfI�?v             g@�       �                    �?(����7�?>            @V@������������������������       �     ��?             @@������������������������       �T�7�s��?*            �L@�       �                    �?�q�Q�?8             X@������������������������       �z�G�z�?             9@������������������������       ��ګH9�?%            �Q@�       �                    �?���Z
�?F           &�@�       �                    �?��W�0��?           ԕ@������������������������       �                     @�       �                    �?T�����?}           ȕ@�       �                     �?�3�c�?�           ��@������������������������       ������Q�?�            �v@������������������������       �����8�?�            �r@�       �                     �?<vhm�B�?�           �@�       �                    �?�Qo�T��?            {@������������������������       ��u����?�             q@������������������������       ��A��4�?_            �c@�       �                    �?�Tޫvɼ?�            �r@������������������������       �`�f��?n            �d@������������������������       �X�Հ�+�?W            �`@�       �                     �?P7�?�           x�@�       �                    �?0G�}i��?h           P�@�       �                    �?�!=�?�           ȇ@������������������������       �0�4ɇ�?>           @������������������������       �X�l�ؾ?�            �p@������������������������       ����K ]�?�             n@�       �                    �?!W[ �?_           ��@������������������������       ����$�?           P{@�       �                    �?�S`1DK�?C           �@������������������������       ��>	<2�?�            �k@������������������������       ��8���?�             r@�       h                   �?�����?/0          �&�@�       E                   �?ʒ�z[��?            �@�       *                   �?�ǫz���?�
           ��@�                          �?�`���?           ��@�                          �?�y�rF�?�           ��@�       �                    �?�s�����?            {@�       �                     �?HP�s��?@             Y@�       �                    �?���N8�?             5@������������������������       �r�q��?             2@������������������������       ��q�q�?             @�       �                    �?(�5�f��?1            �S@������������������������       � ��WV�?0            �S@������������������������       �                     �?�       �                     �?���6���?�            �t@�       �                    �?v�2t5�?k            �d@�       �                    �?�O�y���?a            �b@������������������������       �<W#.m��?E            @Z@������������������������       �z�G�z�?            �F@������������������������       �        
             ,@                          �?0�t�\�?r            @e@                         �?,�Ѡ���?m            �d@������������������������       ��ʻ����?W             a@������������������������       �      �?             <@������������������������       �                     @                         �?u�6/��?�           ,�@                          �?�F��0�?           |�@                         �?�y����?p           ��@������������������������       �                     @	      
                   �?���<_�?m           p�@������������������������       �        l            �f@������������������������       �x�����?           �y@                         �?���N8�?�           X�@������������������������       �                     @                         �?@����u�?�            �@������������������������       ���즟E�?v            �e@������������������������       ����v֧�?           P}@                         �?����z��?{           `�@                          �?@�:;��?o            �f@������������������������       �        B            �[@������������������������       �`����֜?-            �Q@                          �?D�ޢL3�?           p{@������������������������       ��>��(+�?�             o@������������������������       �\�ih�<�?}            �g@                         �?pIC'�T�?           ��@                          �? 7���B�?             ;@������������������������       �                      @������������������������       ��}�+r��?             3@      #                    �?��Oi��?o           �@                          �?LK�?.�?�            �p@                         �?����3��?             J@������������������������       ����X�K�?            �F@������������������������       �؇���X�?             @!      "                   �?�HGݐ\�?�            `k@������������������������       �                    �F@������������������������       ��d���?h            �e@$      '                   �?�}P@�?�             s@%      &                   �?d}h���?/            �Q@������������������������       �     ��?+             P@������������������������       �                     @(      )                   �?_k,D	�?�            �m@������������������������       �(L���?            �E@������������������������       �����ڽ?             h@+      8                    �?@?5�i��?�           ��@,      -                   �?�'֞��?{           ��@������������������������       �                     <@.      3                   �?��Eʸ�?j            �@/      0                   �?`��Ҙ�?�            �t@������������������������       �@f����?l            �c@1      2                   �?��Bs�?g            �e@������������������������       �P����?!            �M@������������������������       �0�)AU��?F            �\@4      7                   �?>�r����?�            �n@5      6                   �? s8TI�?m            �f@������������������������       �FVQ&�?J            �`@������������������������       ��w��#��?#             I@������������������������       ��n_Y�K�?*            @P@9      :                   �?�;�RC�?\           X�@������������������������       �        4            �S@;      @                   �?7�aR=�?(           ��@<      =                   �?`ء�}��?X           ��@������������������������       �@�`%���?�            `r@>      ?                   �?���Ԋ"�?�            `q@������������������������       � ���J��?+            �S@������������������������       ��(\����?x             i@A      D                   �?�z�Ga�?�             t@B      C                   �?nM`����?�            �l@������������������������       �����|-�?q             f@������������������������       ��q�q�?$             K@������������������������       �*;L]n�?;            �V@F      W                   �?t��:���?            �@G      P                   �?�t�&�$�?l           �@H      I                   �?�=����?            z@������������������������       �                     <@J      M                   �?���t��?�            `x@K      L                    �?겡L ��?�            �p@������������������������       ��<<�څ�?S            ``@������������������������       �">�֕�?_            �a@N      O                    �?^;|��?E            �]@������������������������       �"pc�
�?%            �P@������������������������       �H(���o�?             �J@Q      T                    �?~|z����?d            �c@R      S                   �?�5��?%             K@������������������������       �                     "@������������������������       ����X�K�?             �F@U      V                   �?p�9�A��??            @Z@������������������������       �                     4@������������������������       �Ї?��f�?3            @U@X      a                   �?���T�?�           ��@Y      Z                   �?�W�a=�?�           ��@������������������������       �                     $@[      ^                    �?@݈g>h�?�           Б@\      ]                   �?�E���?q           ��@������������������������       ��z�a�?            `y@������������������������       � �Cc}�?q             e@_      `                   �?�����?q           ��@������������������������       �������?            z@������������������������       �HP�s��?a            �b@b      e                    �?��o���?�           �@c      d                   �?0_�n~f�?�            0p@������������������������       �                     @������������������������       ���S�ۿ?�            �o@f      g                   �?�G���?           �{@������������������������       �                     @������������������������       ����*�D�?           �{@i      �                   �?N�u�P��?            ��@j      �                   �?8����?	           ��@k      |                    �?l�+� ��?@           ��@l      w                   �?�~�rR��?            z@m      p                   �? �@*��?�            �q@n      o                   �?l���u�?�            `n@������������������������       ��8��8��?�             k@������������������������       �l��
I��?             ;@q      t                   �?�Gi����?            �B@r      s                   �?��S�ۿ?             .@������������������������       ������H�?             "@������������������������       �                     @u      v                   �?���7�?             6@������������������������       ��X�<ݺ?             2@������������������������       �                     @x      {                   �?�nkK�?T            @a@y      z                   �?�h����?F             \@������������������������       �h㱪��?D            �[@������������������������       �                      @������������������������       �                     :@}      �                   �?�7��d��?:            �@~                         �?�ת2�%�?]           `�@������������������������       �`�0����?8           �~@�      �                   �?��a�n`�?%             O@������������������������       ����|���?             &@������������������������       �`'�J�?            �I@�      �                   �? ~�����?�            �u@�      �                   �?d�
��?             F@������������������������       ��q�q�?             ;@�      �                   �?�t����?             1@������������������������       ������H�?             "@������������������������       �      �?              @�      �                   �? "��u�?�            �r@������������������������       �Pa�	�?�            �p@�      �                   �?�E��ӭ�?             B@������������������������       �                     @������������������������       �ܷ��?��?             =@�      �                    �?,��:��?�           l�@�      �                   �?\���HC�?�           (�@�      �                   �?(�S�,�?�           ȇ@�      �                   �? &;�i�?a           ��@�      �                   �?H����?           0z@������������������������       � ���v�?T             a@������������������������       ��*/�8V�?�            �q@������������������������       ��U���?Q             _@�      �                   �?������?�            @k@������������������������       �@3����?#             K@�      �                   �?�{�����?l            �d@������������������������       ���U�=��?W            �`@������������������������       �      �?             @@�      �                   �?b��L��?�            u@�      �                   �?���؅��?�            �m@������������������������       �p���?             I@������������������������       �d۬����?s            @g@������������������������       ��g��@(�?A            @Y@�      �                   �?�^qj�{�?           ��@�      �                   �?� QG���?3           ��@�      �                   �?��E)���?�           H�@�      �                   �?���a�!�?&           �}@������������������������       �������?U             a@������������������������       � �ʚ�,�?�            u@������������������������       ��zv�X�?u             f@�      �                   �?p3����?�            �m@�      �                   �?\� ���?|            �h@������������������������       �                    �B@������������������������       �0��_��?d            �c@������������������������       �v�2t5�?            �D@�      �                   �?>%Ɍ�S�?�            `w@�      �                   �?|�l�]�?�             q@������������������������       �                      J@������������������������       ��Ra����?�            �k@������������������������       ���.k���?9            �Y@�      �                    �?hh���¼?           ��@�      �                   �?���
�*�?           ĩ@�      �                   �?�)�Z*�?�           (�@�      �                   �?x[�ׂ��?�            �@������������������������       �        T            �@�      �                   �?DGr���?l           @�@������������������������       �ܻ�yX7�?s            @e@������������������������       �����Y�?�           ��@�      �                   �?�ͧ���?�             x@������������������������       �        @             ]@�      �                   �?���"��?�            �p@������������������������       ��q�q�?            �F@������������������������       ����
���?�             l@�      �                   �?�~A���?\           `�@������������������������       ��&6�v�q?!           �|@�      �                   �?(J��_!�?;           P�@������������������������       ��P�*�?P             _@������������������������       ��A5�B�?�           p�@�      �                   �?85Ո醼?           \�@�      �                   �?h+��n��?�           ��@�      �                   �?�K� ��?X           f�@������������������������       �@���?�           8�@�      �                   �?TޓM_�?�           ��@������������������������       �^������?�            �n@������������������������       ��n�Y��?           ��@�      �                   �?x�V�|��?R           8�@�      �                   �?�������?o             g@������������������������       ��6H�Z�?G            @]@������������������������       ��ʻ����?(             Q@������������������������       �8��"s�?�            �v@�      �                   �?�ҵO!�?W           �@������������������������       � �7��p?}           �@�      �                   �?|��8Wv�?�           �@������������������������       ���|�	��?x            �f@������������������������       �����v�?b           <�@rD  trE  bh�h"h#K �rF  h%�rG  RrH  (KM�KK�rI  hQ�B0      �c�@    ���@     ��@     <�@    �[�@     Ԝ@    ��@     <�@      j@     �k@     ��@     ��@     �@     �o@     �y@     �o@     �p@     @n@     `e@     �V@     @W@     �b@     �b@      (@     �_@      &@     �Y@      @     @Y@      @      �?              9@      @      8@      �?      4@              @      �?     �k@            �h�@     ��@    �?�@     �t@     ��@     @Z@     ��@     �H@     (�@     �A@     H�@      @@     Ȁ@      ;@       @             ��@      ;@      q@      @      N@      @      9@      @     �A@              G@      ,@      B@      ,@      $@             �v@      L@     �t@     �K@     �s@      C@     @i@     �A@     �[@      @      4@      1@      =@      �?      1@      �?      (@             ��@     �k@     ��@      .@     ��@       @     ȕ@       @     ,�@             (�@      *@     ��@      *@     ��@             ;�@      j@     ��@     �Y@     (�@      P@     ؄@     �C@     ��@     @Z@     p�@     �S@     ��@     �E@     ��@     �A@     �{@      ;@     �o@      ,@     �g@      *@     ��@     �v@     �r@     `f@     @k@     �U@      i@     �T@      g@      J@     �]@     �B@     �P@      .@      .@      ?@      2@      @      $@       @       @      �?      T@     @W@      �?      �?     �S@      W@      N@     @V@      @@     �M@      <@      >@      3@      .@      "@      .@      3@      @      &@      @      @      �?      @       @       @             P�@      g@     �@      5@     ��@      0@     �v@      $@     �p@      @     H�@      @     x@      @     �m@       @     �b@      �?      a@       @     �U@      �?      I@      �?     ��@     `d@     �@     �T@     @}@     �B@     �t@     �F@     x�@     @T@     @�@     �I@      y@     �@@     �f@      2@     pt@      >@     �m@      8@     �V@      @     `�@     0�@     h�@     u@      @      =@       @      3@              (@       @      @       @       @              @      @      $@      @       @      @      @      �?      �?               @     8�@     @s@     �@     `q@     `v@      c@     �j@      [@      b@     �F@       @             �a@     �F@     �o@     @_@     �a@     �V@     �[@      A@      Y@      >@     �M@      1@     �D@      *@     �|@     Pu@      j@      e@     �[@      Y@              &@     �[@     @V@     @X@      Q@              $@     @X@      M@     `o@     �e@      c@     �X@      Z@     @Q@       @       @     �Y@     �P@      H@      =@              @      H@      7@     �X@     �R@              3@     �X@      L@      P@      >@     �A@      :@     ؂@     �@     �v@     ��@      B@     ��@      2@     `|@      (@     �p@      &@      `@              �?      &@     �_@      �?     �a@      @      g@      @      L@              @@      @      8@       @      `@       @     �F@             �T@      2@     �y@      $@     t@               @      $@     �s@      "@     �n@      @      W@      @      c@      �?     @Q@      �?      ?@              C@       @     �U@      @      C@      @     �H@     pt@     0�@     �p@     0�@     `e@     `t@     �W@      e@      H@      \@     �G@      L@      S@     �c@      J@     �U@      8@      R@     �X@      h@     �O@     @X@      B@     �M@      ;@      C@      B@     �W@      4@     �M@      0@      B@     �L@      `@      A@     �K@      "@      7@      9@      @@      7@     @R@      @      4@      2@     �J@      n@     F�@     ``@     ȓ@              @     ``@     ��@      P@     ��@     �B@     �t@      ;@     �p@     �P@     Є@     �H@     �w@      >@     �n@      3@     `a@      2@     �q@      &@     `c@      @      `@     @[@     Ĝ@      O@     `�@     �D@     ��@      8@     �}@      1@     �n@      5@     �k@     �G@     (�@      1@     @z@      >@     ~@      .@     �i@      .@     0q@     |�@     �@     ��@     f�@     ��@     ��@     �@      ~@     ��@     �u@      f@     p@       @      W@      @      0@      @      .@       @      �?      @      S@      @     �R@              �?      e@     �d@      X@      Q@     �T@      Q@      G@     �M@      B@      "@      ,@             @R@     @X@     �P@     @X@      N@      S@      @      5@      @             Л@     �U@     Ē@      G@     (�@      .@      @             ��@      .@     �f@             �x@      .@     `�@      ?@      @             (�@      ?@     �e@      �?     p{@      >@     �@     �D@     �f@      �?     �[@             @Q@      �?     �x@      D@     `m@      ,@     �d@      :@     @}@      a@      �?      :@               @      �?      2@     0}@     �[@     @m@     �B@      3@     �@@      *@      @@      @      �?     �j@      @     �F@             @e@      @      m@     @R@      .@     �K@      "@     �K@      @             @k@      2@     �B@      @     �f@      (@     �k@     $�@     @V@     �@              <@     @V@     p~@      @     Pt@      �?     `c@      @     @e@      �?      M@       @      \@     @U@     @d@      N@     �^@     �E@     @V@      1@     �@@      9@      D@     �`@     0�@             �S@     �`@     ��@      "@     ��@       @     @r@      @     �p@       @      S@      @     `h@      _@     �h@     @U@      b@     �P@     @[@      2@      B@     �C@     �I@     `@     (�@     `v@     `k@      q@      b@              <@      q@      ]@     @g@     @U@     �V@     �D@      X@      F@      V@      ?@      K@      (@      A@      3@      U@     �R@      @@      6@              "@      @@      *@      J@     �J@              4@      J@     �@@      b@     ��@     @Z@     T�@              $@     @Z@     ,�@     �Q@     p@     �J@     v@      2@     �b@      A@     ��@      6@     �x@      (@     @a@     �C@     Є@      1@     @n@              @      1@     �m@      6@     �z@              @      6@     0z@     ^�@    ���@     (�@      �@     �[@     ��@     �G@     0w@     �D@     �m@      :@      k@      2@     �h@       @      3@      .@      6@      ,@      �?       @      �?      @              �?      5@      �?      1@              @      @     �`@      @     �Z@      @     �Z@       @                      :@     �O@     (�@      8@     ��@      2@     �}@      @      L@      @      @       @     �H@     �C@     s@      5@      7@      "@      2@      (@      @       @      �?      @      @      2@     �q@       @      p@      $@      :@      @              @      :@     ��@      y@     0�@     �d@     h�@      [@     �|@     �T@     0x@      @@     �`@       @     �o@      >@     �R@      I@      h@      :@     �J@      �?     `a@      9@     �\@      1@      8@       @     �q@      L@     �j@      7@     �H@      �?     �d@      6@      Q@     �@@      �@     �m@     Ȇ@     �c@     `�@     @_@      z@     �L@     @_@      &@     0r@      G@      [@      Q@     �i@      @@     �f@      .@     �B@              b@      .@      8@      1@     pr@     �S@     �n@      9@      J@             `h@      9@      H@      K@     ؀@    ���@      i@     4�@      [@     x�@     @U@     ̖@              �@     @U@     ��@      C@     �`@     �G@     x�@      7@     �v@              ]@      7@     �n@      .@      >@       @      k@      W@     �@      �?     �|@     �V@     x�@      J@      R@     �C@     8�@     0u@     	�@     @i@      �@     �b@     8�@      @     $�@     @b@     L�@      U@      d@      O@     Ȓ@     �I@     @@      ?@     @c@      �?      ]@      >@      C@      4@     �u@      a@     �@       @     ؏@     �`@     ��@      O@      ^@     @R@     �@rJ  trK  bubhhubh)�rL  }rM  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h7Kh8Kh9h"h#K �rN  h%�rO  RrP  (KK�rQ  hQ�C              �?rR  trS  bhEhUh@C       rT  �rU  RrV  hYKhZh[Kh"h#K �rW  h%�rX  RrY  (KK�rZ  h@�C       r[  tr\  bK�r]  Rr^  }r_  (hKheM�hfh"h#K �r`  h%�ra  Rrb  (KM��rc  hm�Bc         2                   �?��A2��?�e           �@       �                     �?��B+��?�9          @��@       j                    �?�q�����?*"          ��@       	                    �?xaE�Q�?�          ���@                           �?�c���?�           ��@                            �?flx����?�           ��@������������������������       ���*��?           �{@������������������������       ��
X���?�            `o@������������������������       �                     @
       5                    �?\3 0��?D          �\�@       $                    �?�'N��?�           ��@                           �?({��i�?U           ܔ@                           �?�hrF��?           p�@                           �?��7N�?�           X�@                           �?P>�F�?\           ��@                           �?�Q�9�ϱ?�           Ȅ@������������������������       ��q�q�?=             X@������������������������       ��Un� ܳ?c           ȁ@                           �?PpS�Ж�?�            �q@������������������������       �                     (@������������������������       ��(�T[X�?�             q@                           �?R۔t��?�            �k@������������������������       ���+7��?]            @a@������������������������       ��ucQ?-�?6            @U@                           �?`����֜?+            �Q@                           �?�h����?#             L@                           �?�nkK�?             7@������������������������       �                     �?������������������������       ����7�?             6@������������������������       �                    �@@������������������������       �                     ,@        #                    �?��|�	��?;            �V@!       "                    �?l�;�	�?1            �R@������������������������       ���+7��?             G@������������������������       �J�8���?             =@������������������������       �        
             0@%       4                    �?�z�X���?�           H�@&       /                    �?�\��9�?k           ��@'       ,                    �?�Y�R_�?           �z@(       +                    �?|6����?�             u@)       *                    �?     ��?S             `@������������������������       ��q�q�?             B@������������������������       �\X��t�??             W@������������������������       �\�����?�            @j@-       .                    �?�0�~�4�?5             V@������������������������       �F�t�K��?             �L@������������������������       �f���M�?             ?@0       3                    �?<���|��?\            @a@1       2                    �?��k=.��?            �G@������������������������       �                      @������������������������       ��θ�?            �C@������������������������       �p�C��?=            �V@������������������������       �                    �J@6       S                    �?���?e          ���@7       H                    �?����&"�?�           ׺@8       A                    �?����t�?=           ��@9       >                    �?�qI��5|?"           ��@:       =                    �?���Lj�q?�           J�@;       <                    �?���H��?�           t�@������������������������       �        B            @[@������������������������       � *t:#l�?U           ��@������������������������       �        &            �@?       @                    �?��˼��?e             e@������������������������       �                     @������������������������       �������?a            `d@B       C                    �?�I�Z�?           ��@������������������������       �                     @D       G                    �?8օ{�d�?           ��@E       F                    �? �}FQ�?]           <�@������������������������       ����&B�?�           \�@������������������������       � "�4 ڮ?i           �@������������������������       �`�dG�?�            �r@I       N                    �?P~�2�,�?�           ��@J       K                    �?@ѽ�֞?�            pt@������������������������       �                     "@L       M                    �?`I�)豟?�            �s@������������������������       �����?r             f@������������������������       �        \            �a@O       P                    �?�J�lc+�?�           ��@������������������������       ��kb97�?�            x@Q       R                    �?���.�6�?�             w@������������������������       �x�U���?�            �m@������������������������       � �#�Ѵ�?W             `@T       _                    �?йJ	˸?t           ��@U       \                    �? d�ٟ?<           ��@V       Y                    �? ��o� �?�           ��@W       X                    �? _�@�Y�?%            }@������������������������       ����͡?�            0u@������������������������       �@�n�1�?T            @_@Z       [                    �? �.�?Ƞ?�            �r@������������������������       �0��kS֣?�            �o@������������������������       �                    �G@]       ^                    �? ��7��?K            �^@������������������������       �����ȫ�?3            �T@������������������������       �                     D@`       c                    �? 	��p�?8           0�@a       b                    �?��
b��?�           �@������������������������       �P5f7���?)           �}@������������������������       �ףp=
�?�             r@d       g                    �?௩�F��?Z           x�@e       f                    �?8�a$��?|           �@������������������������       ����[�?            �|@������������������������       �Х-��ٹ?\            �b@h       i                    �?��GEI_�?�            �v@������������������������       ��@�?h            `d@������������������������       ����"F��?v            `i@k       x                    �?U�ǲ��?8           �@l       q                    �?Z[��-O�?           `�@m       n                    �?�?�H\�?7           �@������������������������       �                     8@o       p                    �?���,���?*           0~@������������������������       �V�#y��?�             w@������������������������       ��"'`�]�?J            @\@r       u                    �?������?�            u@s       t                    �?�חF�P�?             ?@������������������������       �ףp=
�?             $@������������������������       ���s����?             5@v       w                    �?�zܯ�V�?�             s@������������������������       ��	��c��?|             h@������������������������       �VcYE�?H            @\@y       �                    �?6P�����?(           p�@z                           �?��\���?W            �@{       ~                    �?�J�4�?             9@|       }                    �?����X�?	             ,@������������������������       ����!pc�?             &@������������������������       ��q�q�?             @������������������������       �                     &@�       �                    �?BH7�B�?G           8�@�       �                    �?���B���?            z@������������������������       ��"U����?�            �o@������������������������       �pa�M���?e             d@�       �                    �?�O��i�?A            �Y@������������������������       ��z�G��?'             N@������������������������       ���V#�?            �E@�       �                    �?�k���)�?�            �t@�       �                    �?��(\���?             D@�       �                    �?P���Q�?             4@������������������������       �؇���X�?             @������������������������       �                     *@�       �                    �?ףp=
�?             4@������������������������       �                     @������������������������       ��t����?             1@�       �                    �?��tT"�?�            `r@�       �                    �?=��T�?Y            �a@������������������������       ���V#�?             �E@������������������������       ���ga�?9            @X@�       �                    �?�X����?_            @c@������������������������       �     ��?&             P@������������������������       �F�����?9            �V@�       �                    �?P�D�~�?�           ��@�       �                    �?������?�           \�@�       �                    �?�p0`���?�           d�@�       �                    �?d:���?�             w@�       �                    �?�j4/��?�            pp@�       �                    �?�wh�?�            p@������������������������       ��k�ɲ��?�             m@������������������������       ��q�q�?             8@������������������������       �r�q��?             @�       �                    �?P�c0"�?F            @Z@������������������������       �F|/ߨ�?7            @T@������������������������       �                     8@�       �                    �?�T/�rZ�?�           H�@�       �                    �?b*ꃮ��?�           �@�       �                    �?�ӭ�a��?            {@�       �                    �?��z��1�?�            �x@������������������������       �                      @�       �                    �?�X�C�?�            �x@�       �                    �?�mqA{��?�            �u@������������������������       �2m7a��?�            �l@������������������������       ��1e�3��?M            �]@������������������������       ��q�q�?            �F@�       �                    �?�˹�m��?             C@������������������������       �     ��?	             0@������������������������       �                     6@�       �                    �?��c����?�             q@�       �                    �?�<,Ҫ��?�            �i@�       �                    �?V��f_�?|            �h@������������������������       ��G�z��?b             d@������������������������       �      �?             B@������������������������       �                     "@�       �                    �? ���g=�?+            @Q@������������������������       ��i�y�?'            �O@������������������������       �                     @�       �                    �?�θ�?            �C@�       �                    �?�z�G��?             >@�       �                    �?8����?             7@������������������������       ����|���?             &@������������������������       �      �?             (@�       �                    �?����X�?             @������������������������       �      �?             @������������������������       �                     @������������������������       �                     "@�       �                    �?��nm���?�           T�@�       �                    �?fn�
>�?�           x�@�       �                    �?@u��?�           8�@�       �                    �?�Ƀ aA�?H            �]@������������������������       ��q�q�?             @�       �                    �?��|��L�?E            �\@�       �                    �?�/���??            �Y@������������������������       ���c:�?9             W@������������������������       �                     &@������������������������       �                     (@�       �                    �?�IFz�?O           ��@������������������������       ���j:|�?+           �}@�       �                    �?H%u��?$             I@������������������������       ��q�q�?             @������������������������       ����7�?              F@�       �                    �?$��m��?@             Z@�       �                    �?(����7�?6            @V@�       �                    �?`�Q��?.            �R@������������������������       ��4�����?             ?@������������������������       �t��ճC�?             F@�       �                    �?����X�?             ,@������������������������       �      �?              @������������������������       ��q�q�?             @�       �                    �?�r����?
             .@������������������������       �                     "@������������������������       ��q�q�?             @�       �                    �?p�լ�?�?�            `v@�       �                    �?(�T����?�            �r@������������������������       �V�a�� �?             =@������������������������       ���}����?�            �p@�       �                    �?`��:�?(            �N@�       �                    �?$�q-�?             *@������������������������       �                     @������������������������       ������H�?             "@������������������������       �                     H@�                          �?ІW#�N�?@           ̼@�                          �?�eP-Q�?�           ��@�       �                    �?�G�N�*�?�	           Ю@�       �                    �?������?>           ܙ@������������������������       �                     E@�       �                    �? �g�s_�?'           4�@�       �                    �?��G^�C�?           H�@�       �                    �? �jY6;�?�           ��@������������������������       ���r6��?�           8�@������������������������       �        1           p}@������������������������       ��Ń��̧?;             U@�       �                    �? �ؒ;S�?"           �{@������������������������       �@Lb�G�?�            @o@�       �                    �? bB���?~             h@������������������������       �@�`%���?a            `b@������������������������       �                     G@�       �                    �?�Q�E�(�?�           �@�       �                    �?��y��?�           �@�       �                    �?�4{r�ٸ?b           ��@�       �                    �?0�ج �?�           h�@������������������������       �                     @������������������������       �`��X�?�           0�@�       �                    �?�k3����?�           ��@������������������������       �                     @������������������������       �H�*�ɺ?�           ��@������������������������       �$Nz�{�?�             k@�                          �?$l�q[��?�           `�@�                           �?����?i           ��@������������������������       �ףp=
�?�             t@������������������������       ���O���?�            �o@������������������������       � '��h�?B            @[@      
                   �?��?��?           0�@                         �?     G�?�            �@                         �?�+��b�?U           �@������������������������       �p�`Bh�?g            �b@������������������������       �K����?�            �x@      	                   �?���R���?+           �}@������������������������       � �q�q�?P             ^@������������������������       �H�73m��?�            Pv@                         �?�p�O�A�?�           `�@                         �?��8�$>�?~            @h@                         �?��s�n�?C             Z@                         �?F��}��?2            @R@������������������������       �                     �?������������������������       ��X�<ݺ?1             R@������������������������       ��g�y��?             ?@                         �?(;L]n�?;            �V@������������������������       ���(\���?             D@������������������������       �        !             I@                         �?�`it)�?           ��@                         �?`���i��?           �{@������������������������       ��e)���?�            �m@������������������������       ����"F��?�            `i@                         �?���>W�?�            �y@������������������������       �h��@D��?Y            �a@������������������������       �l��\��?�             q@      '                   �?v�!��?b           0�@      "                   �?�+v���?�           ��@                         �?P;8����?           �y@������������������������       �Ȩ�I��?�            �j@       !                   �?���!x��?�            @i@������������������������       �~�u���?[            �a@������������������������       ���Q:��?'            �M@#      $                   �?RŪx���?�            ps@������������������������       ��J�T�?[            �a@%      &                   �?nmR���?m             e@������������������������       ��\��N��?=            �W@������������������������       �      �?0            �R@(      -                   �?��697�?�           ��@)      *                   �?θ	j*�?�            �s@������������������������       ��T���?^            `d@+      ,                   �?��s��?]            �b@������������������������       �rr�J��?(            �R@������������������������       ���H�}�?5            �R@.      1                   �?�*n�x�?�            �s@/      0                   �?2e�3���?�            �m@������������������������       �0S>�U�?s            �f@������������������������       �      �?$             L@������������������������       �|jq��?:            �T@3      |                   �?:{�~�?�+          �P�@4      c                   �?��/�g��?�           <�@5      L                   �?(i�qْ�?�           t�@6      A                   �?�GN�z�?G           0�@7      >                   �?8��H��?            y@8      =                   �?X]�hx�?�            ps@9      :                   �?xsG��?�             m@������������������������       �                     @;      <                    �?�D�n���?�            `l@������������������������       ����.�d�?^            �a@������������������������       ��D�e���??            @U@������������������������       �        5            �S@?      @                    �?4�<����?6            @V@������������������������       �:	��ʵ�?            �F@������������������������       ��C��2(�?             F@B      I                   �?:�6���?:           `@C      F                    �?f������?           0z@D      E                   �?P&��?�            �m@������������������������       ��S��<�?Y            �a@������������������������       �0d4�[%�?;            �W@G      H                   �?����W��?s            �f@������������������������       ��q�q�?D            �X@������������������������       ��i#[��?/             U@J      K                    �?NP�<��?3            �T@������������������������       �H.�!���?             I@������������������������       ��eP*L��?            �@@M      X                   �?�޶��?p           ��@N      U                   �? w���%�?h           ��@O      R                    �?@�-	�?           pz@P      Q                   �?�K��h�?�            �h@������������������������       � E��ۛ?^             b@������������������������       �@3����?#             K@S      T                   �?����X�?�             l@������������������������       ��E�����?k            �f@������������������������       �                     F@V      W                    �? i�*$Ŋ?`             c@������������������������       � }�Я��?8            @V@������������������������       �        (            �O@Y      `                   �?ȐY"��?           �y@Z      ]                    �?����X�?�            @s@[      \                   �?�1��n�?w            �e@������������������������       �4և��P�?M             \@������������������������       �Nd^����?*            �N@^      _                   �?L/)Lr��?X            �`@������������������������       �>��C��?;            �U@������������������������       ��q��/��?            �H@a      b                    �?��:M�?9             Y@������������������������       ��99lMt�?            �C@������������������������       ��ɞ`s�?            �N@d      o                    �?� O��?0           ��@e      j                   �?(�P���?N           @�@f      i                   �?�A�D6h�?           �@g      h                   �?@݈g>h�?�           `�@������������������������       ���y/���?           �y@������������������������       �0M����?�            �p@������������������������       �̻L&��?Y            �b@k      l                   �?m��"2�?L           h�@������������������������       ���92��?           �{@m      n                   �?(�1uԳ�?.           �|@������������������������       �`�I��g�?�            �l@������������������������       ��8h
Q��?�             m@p      w                   �?�I &���?�           <�@q      r                   �?L:�f@�?�           ��@������������������������       �                      @s      t                   �?\���R�?�           Ђ@������������������������       ��:pΈ��?�            �r@u      v                   �?@�+9\J�?�            �r@������������������������       �����\�?r            �f@������������������������       ���GEI_�?O            �^@x      {                   �?pN�{Mb�?]           ��@y      z                   �?�04��X�?�           ��@������������������������       ���z�}�?           �{@������������������������       ��*E
S�?�            �l@������������������������       �@��9U��?�            @q@}      �                   �?�L)�2�?�          ���@~                         �?�������?�           *�@������������������������       �        [            �`@�      �                   �?$2#po��?)           �@�      �                   �? ���`�?M           �@�      �                   �?4)�ʀ�?           4�@�      �                    �?�!����?.           p~@������������������������       ��f]/U�?v            �g@������������������������       � c�O�?�            �r@�      �                   �?n)�z8��?�           ��@�      �                    �?�<�.W�?�            �r@������������������������       �VcYE�?I            @\@������������������������       �x������?|            �g@�      �                    �?$H/E��?           ��@������������������������       �H��3rY�?�            �w@������������������������       ��Պ&�4�?           �{@�      �                    �?0a�G�?J           X�@�      �                   �?V�g�8~�?�            `o@������������������������       ���?^�k�?            �A@�      �                   �?�+$�jP�?}             k@������������������������       ��&�5y�?!             O@������������������������       �vl��C�?\            @c@�      �                   �?��)�c{�?�             s@������������������������       ���+��<�?,            �U@�      �                   �?�A�m��?�            @k@������������������������       ����Q��?              I@������������������������       �l������?j             e@�      �                   �?</z���?�           X�@�      �                    �?�����?           |@�      �                   �?�+$�jP�?w             k@������������������������       ��U���?F            �_@������������������������       �ƈ�VM�?1            @V@�      �                   �?����?�             m@������������������������       �@�E�x�?f            `b@������������������������       �t���D�?:            �U@�      �                    �? )�y���?�           ��@������������������������       ��Q�p6м?�            �q@������������������������       �X�QnO�?           �{@�      �                    �?��,��?T           ��@�      �                   �?�:��h`�??           ��@�      �                   �?�\1�K3v?�           @�@�      �                   �? .���4i?�           H�@������������������������       � L�C��n?b           ��@������������������������       �        ?            @\@������������������������       � [ĉ��?$           p|@�      �                   �?�J��Ed�?z           X�@�      �                   �?l�X�e�?            �@������������������������       ��
���K�?o            �e@������������������������       ��j�$�e�?           ؊@�      �                   �?W�!?�?�           ��@�      �                   �?�A��4�?�            �s@������������������������       ��n_Y�K�?!            @P@������������������������       ���H�$�?�            `o@�      �                   �?xE(�B��?7           @�@������������������������       �V{q֛w�?S             _@������������������������       �+Rh�r�?�           `�@�      �                   �?p���1�?           v�@�      �                   �? ~���?�           ҡ@������������������������       � '�vf�}?�           4�@�      �                   �?�� �JH�?�           p�@������������������������       ��P[1N�?^            �b@������������������������       � FR2Ш?�           �@�      �                   �?�ox��X�?           �@�      �                   �?�q�q�?]           X�@�      �                   �?�2�2�?�             u@������������������������       ���T�l��?�            �p@������������������������       ���%��?+            �R@������������������������       �>����?�             k@�      �                   �?�X;�^��?"           Ħ@������������������������       �x��:߷?�           |�@�      �                   �?hG�3;۰?/           �@������������������������       ��l��6�?�             u@������������������������       ��7zD��?\           ̕@rd  tre  bh�h"h#K �rf  h%�rg  Rrh  (KM�KK�ri  hQ�BP       P�@     ��@     ��@     U�@     u�@     �@    �n�@     P�@     pw@     t@      w@     t@     �j@     �l@     �c@     @W@      @             ��@     ��@      �@      �@     �@     �^@      �@      W@     �@     �V@     Ќ@      =@     �@      8@     �W@      �?     �@      7@     �q@      @      (@             �p@      @      d@      O@     �Y@      B@     �M@      :@     @Q@      �?     �K@      �?      6@      �?      �?              5@      �?     �@@              ,@              N@      ?@      F@      ?@      A@      (@      $@      3@      0@             �h@     Pz@     �a@     Pz@     �`@     `r@     �R@     pp@      J@      S@      (@      8@      D@      J@      7@     `g@     �L@      ?@      G@      &@      &@      4@      &@     �_@      "@      C@               @      "@      >@       @     @V@     �J@             ��@     0s@     *�@     �e@     #�@      _@     ��@      $@     >�@      @     \�@      @     @[@             ��@      @      �@             �d@      @      @             �c@      @     ��@     �\@      @             ��@     �\@     ~�@     �W@     ��@     �I@     l�@      F@     �q@      3@     �@     �H@      t@      @      "@             �s@      @     �e@      @     �a@             (�@      F@     �v@      4@     �u@      8@     �k@      2@     �^@      @     x�@     �`@     @�@      ,@     x�@      *@     �|@       @     �t@      @     �^@       @     pr@      @      o@      @     �G@             @^@      �?     @T@      �?      D@             P�@      ^@     ��@      O@     �{@     �@@     Pp@      =@     ��@      M@     ��@      A@     {@      :@     �a@       @     `u@      8@     `c@       @     `g@      0@     4�@     h�@     8�@     Pt@     0u@      e@              8@     0u@      b@     Pp@     @[@     �S@     �A@     �f@     �c@      @      :@      �?      "@      @      1@     �e@     ``@     �Y@     �V@     @R@      D@     0�@     �v@     @t@     �k@      @      5@      @      $@      @       @      �?       @              &@      t@     �h@      o@     �d@      d@     �W@     @V@      R@     �Q@      @@      E@      2@      =@      ,@     @h@     �a@      @     �B@      �?      3@      �?      @              *@       @      2@              @       @      .@     �g@     �Y@     �U@      K@      =@      ,@     �L@      D@     @Z@     �H@     �H@      .@      L@      A@     f�@     (�@     p�@     ��@     ��@     Ѐ@     �]@     @o@      ]@     `b@     �[@     @b@      W@     �a@      3@      @      @      �?       @     �Y@       @     �S@              8@     �|@      r@      |@      p@     �v@     �P@     �t@     �O@       @             �t@     �O@     �r@      H@     �g@     �D@     �[@      @      >@      .@     �A@      @      *@      @      6@             �T@      h@     �R@     ``@     @P@     ``@     �G@     @\@      2@      2@      "@               @     �N@       @     �N@      @              "@      >@      "@      5@      @      0@      @      @      @      "@       @      @       @       @              @              "@     �a@     0�@      \@     ��@      S@     ؁@      I@      Q@      �?       @     �H@     �P@     �H@      K@      C@      K@      &@                      (@      :@     p@      4@     �|@      @      F@      @       @       @      E@      B@      Q@      A@     �K@      8@     �I@      5@      $@      @     �D@      $@      @      @       @      @       @       @      *@              "@       @      @      ?@     pt@      3@     `q@      @      7@      *@     �o@      (@     �H@      (@      �?      @               @      �?              H@     ��@     ��@     9�@     pt@     ��@     @d@     ��@      *@      E@              �@      *@     $�@      "@     ܐ@      @      �@      @     p}@             �T@       @     p{@      @     �n@      @      h@      �?     @b@      �?      G@             ��@     �b@     ��@      V@     ��@     �Q@     X�@      A@      @              �@      A@     Ѓ@     �B@      @             ��@     �B@      i@      1@     x�@     �N@     8�@      L@      r@      @@     �l@      8@      Z@      @     ̝@     �d@     `�@      U@     @�@      ;@     `b@      @     Pw@      7@     @z@     �L@     �\@      @     s@      J@     8�@     @T@     @g@       @     �X@      @     @Q@      @      �?              Q@      @      >@      �?     �U@      @     �B@      @      I@             h�@     @R@     Py@     �A@     @k@      3@     `g@      0@     �w@      C@      `@      ,@      o@      8@     ��@     �~@     �}@     �o@      r@      _@     �c@      L@     �`@      Q@     @X@      G@     �B@      6@     �f@      `@      X@      G@     �U@     �T@      I@     �F@     �B@     �B@     `x@      n@     @j@     �Y@     @]@      G@     @W@      L@     �F@      =@      H@      ;@     �f@     `a@     ``@     @Z@     �Y@     @S@      <@      <@     �H@      A@     ��@    ���@     �@     ٱ@     �t@     D�@     �i@     ȅ@      7@     �w@      &@     �r@      &@     �k@              @      &@      k@      "@     �`@       @     �T@             �S@      (@     @S@       @     �B@      @      D@     �f@      t@     �c@     pp@     �T@     @c@     �J@      V@      =@     �P@     �R@     @[@     �@@     �P@     �D@     �E@      :@     �L@      &@     �C@      .@      2@     �_@     ��@      @     ȁ@      @      z@      @     �h@       @     �a@      �?     �J@       @     �k@       @     @f@              F@      �?     �b@      �?      V@             �O@     @^@     �q@      V@     �k@      O@     �[@     �B@     �R@      9@      B@      :@     @[@      4@     �P@      @     �E@     �@@     �P@      ,@      9@      3@      E@     pq@     ��@     `c@     Ԙ@     @U@     p�@     �O@     h�@     �E@      w@      4@     `o@      6@      `@     �Q@     8�@      =@      z@     �D@     Pz@      4@      j@      5@     �j@      _@     L�@      P@     ��@               @      P@     Ѐ@      E@      p@      6@     �q@      ,@     �d@       @     �\@      N@     ��@      G@     ��@      ;@     �y@      3@     �j@      ,@     `p@     h�@     ��@     �w@     2�@             �`@     �w@     $�@     �p@     ��@     �f@     `�@      @     ~@      �?     �g@      @     0r@     �e@     ��@     @]@     @g@      D@     @R@     @S@     @\@      M@     �@     �@@     �u@      9@     0z@     �T@     �}@     �D@     @j@      �?      A@      D@      f@      1@     �F@      7@     ``@      E@     `p@      @     �T@     �C@     `f@      4@      >@      3@     �b@      ]@     ��@      S@     Pw@      D@      f@      @      _@     �B@      J@      B@     �h@      @      b@     �@@     �J@      D@     h�@      1@     �p@      7@      z@     ��@    ���@     @k@     D�@      @     4�@      �?     @�@      �?     ��@             @\@       @     P|@     �j@     T�@     �W@     H�@      @@     �a@     �O@     ��@      ^@     ��@      C@     `q@      9@      D@      *@     �m@     �T@     ��@      K@     �Q@      <@     ��@     ps@     ?�@      "@     ��@      @     $�@      @     \�@      �?     �b@      @     �@     �r@     ��@      g@      w@     �]@     `k@     @U@     `f@      A@      D@     �P@     �b@     @]@     ڥ@      M@     ��@     �M@      �@      &@     Pt@      H@     �@rj  trk  bubhhubh)�rl  }rm  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h7Kh8Kh9h"h#K �rn  h%�ro  Rrp  (KK�rq  hQ�C              �?rr  trs  bhEhUh@C       rt  �ru  Rrv  hYKhZh[Kh"h#K �rw  h%�rx  Rry  (KK�rz  h@�C       r{  tr|  bK�r}  Rr~  }r  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�B�j         �                    �?���C��?{e           �@       �                    �?�?����?�5           �@                           �?d°�.
�?T(          ���@       	                     �?*�����?g           ��@                            �?
l5p���?�           h�@������������������������       �D���h��?           `|@                           �?�tx>�U�?�            pp@������������������������       ��q�q�?�            Pp@������������������������       �                      @
                           �?��`.��?�            pp@������������������������       ��7�֥��?�            @p@������������������������       �                     @       d                    �?��ʳJ�?�%          ���@       7                    �?�9y��%�?}          �j�@       "                     �?�`Va�?�           x�@                           �?PX����?�           $�@                           �?�nkK�?�           ��@                           �?�}�+K̶?d           p�@                           �?@O��F��?E           �@                           �? >��@�?I            @_@������������������������       � �O�H�?>            �[@������������������������       �                     ,@                           �?x������?�           (�@������������������������       ���+
S,�?N           �@������������������������       �Pns��ޭ?�            �p@                           �?���!pc�?             F@������������������������       �                     �?������������������������       ��%^�?            �E@������������������������       �        (            �Q@       !                    �?؇���X�?             5@                            �?�S����?             3@������������������������       �؇���X�?	             ,@������������������������       �z�G�z�?             @������������������������       �                      @#       (                    �?^�����?.           P}@$       '                    �?     ��?             @@%       &                    �?PN��T'�?             ;@������������������������       ��J�4�?             9@������������������������       �                      @������������������������       �z�G�z�?             @)       2                    �?L��o& �?           P{@*       /                    �?ȵHPS!�?
            z@+       .                    �?�i����?�            Px@,       -                    �?�#c���?�            w@������������������������       �     ��?�             p@������������������������       ��/�z{�?K            @\@������������������������       �                     4@0       1                    �?l��
I��?             ;@������������������������       ��q�q�?             8@������������������������       �                     @3       6                    �?���N8�?             5@4       5                    �?�E��ӭ�?
             2@������������������������       �����X�?             ,@������������������������       �      �?             @������������������������       �                     @8       M                     �?�hto�?�          �{�@9       @                    �?���?�           M�@:       ;                    �? m1�]��?P           ̦@������������������������       �        ?            �X@<       ?                    �?���n�?           �@=       >                    �?��<p��?A           ��@������������������������       �@Wҷ�w�?]           Ԕ@������������������������       ��@)�<�?�           ,�@������������������������       �0�{�F��?�            @t@A       B                    �?8����?^           Ω@������������������������       �        !            �G@C       J                    �?���
1�?=           p�@D       G                    �?�3�R�T�?l           �@E       F                    �? M.[ظ�?E           H�@������������������������       �        �           L�@������������������������       ����?H           D�@H       I                    �?Pl0�ͤ?'            ~@������������������������       �        n             f@������������������������       ��]0��<�?�            s@K       L                    �?�x_F-�?�             s@������������������������       �v�`����?�            @n@������������������������       �     8�?*             P@N       ]                    �?��d5�0�?           T�@O       V                    �?М���}�?             �@P       Q                    �?����?           8�@������������������������       �                    �@@R       U                    �?�Ր�m�?�           ��@S       T                    �?��ht�Y�?�           \�@������������������������       ��g���V�?�           P�@������������������������       ���O�:�p?2           �~@������������������������       ���f�{��?:            �U@W       X                    �?�;Y�&��?�           �@������������������������       �                     $@Y       Z                    �?ʂx���?�           ��@������������������������       ���(��?�           Ȇ@[       \                    �?8��Cu`�?%           ��@������������������������       ��/G�v�?�           (�@������������������������       �H��2�?x            @g@^       a                    �?~j�$s�?           �y@_       `                    �? s�n_Y�?�             j@������������������������       �                     �?������������������������       ��(K\�l�?�            �i@b       c                    �?�#+�f��?�            @i@������������������������       �f�Sc��?^            `b@������������������������       ��b��[��?"            �K@e       �                    �?2��da��?p
           p�@f       w                     �?    �-�?O            �@g       r                    �?R���3�?�            �r@h       m                    �?�� ���?�            �p@i       l                    �?�5�<
�?�            �o@j       k                    �?(�~	WC�?�            �k@������������������������       ���O�;��?W             `@������������������������       ���!���?7            @W@������������������������       �      �?             @@n       q                    �?������?             1@o       p                    �?������?	             .@������������������������       �����X�?             @������������������������       �      �?              @������������������������       �                      @s       t                    �?r�q��?             >@������������������������       �        	             (@u       v                    �?�E��ӭ�?
             2@������������������������       �      �?             $@������������������������       �                      @x       �                    �?:K�����?�            `j@y       �                    �?̕8g���?r             e@z       }                    �?>U���?e            �b@{       |                    �?V�W?�?[             a@������������������������       ����ջ��?A             Z@������������������������       �r٣����?            �@@~                           �?�	j*D�?
             *@������������������������       ��q�q�?             @������������������������       �����X�?             @������������������������       �                     3@�       �                    �?��i#[�?             E@�       �                    �?*O���?             B@������������������������       ��������?             >@������������������������       �                     @������������������������       �                     @�       �                    �?�D��g<�?!	           �@�       �                     �?�N����?A           �@�       �                    �?�d4���?i           �@�       �                    �? ��>��?�           �@������������������������       �`��Ҙ�?�            �t@�       �                    �?�#��Y�u?�            @w@������������������������       �        �             r@������������������������       � ��N8�?1             U@�       �                    �?�t�D��?�           �@������������������������       �X{����?"            ~@�       �                    �?Lea�Y �?�            �@������������������������       �ȴ�S뭽?!           P{@������������������������       �HP�s��?m            �e@�       �                    �?aoMς�?�           Б@�       �                    �? ��fί�?�           �@������������������������       � D�R��?�            q@������������������������       ��l��6�?�             u@�       �                    �?Е�#v��?N           ��@�       �                    �? J���#�?x             f@������������������������       �        V             ^@������������������������       ��h����?"             L@�       �                    �?$'�#�?�            0v@������������������������       �@4և���?�            �o@������������������������       �p�eU}�?B            �Y@�       �                    �?|?n?�?�           ȇ@�       �                    �?�n�q�Z�?�           `�@�       �                     �?�k)Y���?�            Pw@������������������������       �HuWP�x�?�            �j@������������������������       �Z}.�|�?b            �c@�       �                     �?�������?�            �n@������������������������       ��W����?f            �d@������������������������       �F~��7�?:            �T@�       �                     �?ص���?X            �a@������������������������       �*O���?,             R@������������������������       ��q�q�?,            @Q@�       �                    �?l�uwn��?Q           �@�       �                     �?\[�����?�           |�@�       �                    �?h�3��2�?�           Ė@�       �                    �?�ћqQ�?�           ��@�       �                    �?�v��\�?�             q@������������������������       �                     �?�       �                    �?jK�?�j�?�            q@������������������������       ���sK�z�?I            �^@������������������������       ��w��#��?]            �b@������������������������       �Xd,t�?           `z@�       �                    �?h.�Lp�?�           ȇ@�       �                    �?>a�����?�            �o@������������������������       � �kakd�?d            �b@������������������������       �҆�s��?E             Z@������������������������       ����7�?G           �@�       �                    �?�NG�9��?           4�@�       �                    �?*Y�_[�?]           x�@������������������������       �                     "@�       �                    �?�.�	ݗ�?V           0�@������������������������       �h�a��?@            @X@�       �                    �?��o1T��?           P|@������������������������       ����Q��?I             ^@������������������������       �$D�9[�?�            �t@�       �                    �?TKc`�?�           ��@������������������������       ����E�?i            �e@�       �                    �?�Q1t4�?X           ��@������������������������       ��O��i�??            �Y@������������������������       �(M6�tg�?           �|@�       �                    �?�"�a��?�           ��@�       �                    �?��v����?�           �@�       �                     �?�pA��?�           ؆@�       �                    �?���Վ�?           {@�       �                    �?"�����?]            �b@������������������������       �                    �A@������������������������       ���h!��?E            �\@������������������������       �h��@D��?�            �q@�       �                    �?u�����?�            �r@�       �                    �?�q����?C            �Z@������������������������       �                      @�       �                    �?�	j*D�?B             Z@������������������������       ����N8�?             E@������������������������       ��g�y��?&             O@������������������������       ���8����?y             h@�       �                    �?������?�           8�@�       �                     �?@��,B�?<            �V@������������������������       �`���i��?             F@������������������������       �                    �G@�       �                    �?�TL��p�?�           `�@�       �                     �?�������?W            �a@������������������������       ��w���?3            @T@������������������������       �t�7��?$             O@�       �                     �?��:�r�??           �@������������������������       ���W[�?�            �p@������������������������       ��R����?�            @n@�       �                    �?m����?�           L�@�       �                     �?��	2��?�            x@�       �                    �?2H�'�?            �g@�       �                    �?`K�����?0            @R@������������������������       �     ��?             @@������������������������       ��4F����?            �D@�       �                    �?����?O             ]@������������������������       �0�z��?�?+             O@������������������������       ��q�q�?$             K@�       �                    �?ZՏ�m|�?|            �h@�       �                    �?��9J���?B             Z@������������������������       � �#�Ѵ�?            �E@������������������������       ���v$���?'            �N@�       �                    �?�)
;&��?:             W@������������������������       ��E��ӭ�?             B@������������������������       �������?#             L@�       �                     �?���I���?           ��@�       �                    �?h�^����?�            pv@������������������������       ��&1R)�?]            �a@������������������������       �,��J�H�?�            @k@�       �                    �?�-�0�?           �z@�       �                    �?`�BX�l�?Z             a@������������������������       �                      @������������������������       ���S�ۿ?Y            �`@������������������������       � �$@�?�             r@�       ~                   �? .e���?�/           /�@�       U                   �?�Y�)���?�           ;�@�                          �?��=|��?           e�@�                          �?������?�            �k@�                           �?T���.�?�             k@�                          �?�&�5y�?&             O@�                          �?)O���?             B@                          �?l��
I��?             ;@������������������������       � �o_��?             9@������������������������       �      �?              @������������������������       �                     "@������������������������       �                     :@                         �?x�Y��?_            `c@      	                   �?������?:            @V@                         �? 	��p�?8            �U@������������������������       �h�����?6             U@������������������������       �                     @
                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        %            �P@������������������������       �                     @      2                   �?.�&�1��?z           ��@      !                    �?{0����?'           
�@                         �?�T����?�           ��@                         �?��{���?~           �@                         �?�<@�'�?�           ��@                         �?��Q:��?J            �]@������������������������       ��~8�e�?@            �Y@������������������������       �        
             0@                         �?��Ε�X�?x           ؂@������������������������       ��M�a�[�?u            �f@������������������������       � $��*�?           Pz@                         �?��T��g�?�            @s@������������������������       �        o            �f@������������������������       ����Q��?M            @_@                          �?���<�l�?9           ~@                         �?r�����?K            �\@������������������������       �      �?              @������������������������       ���ɜ|��?G            �Z@������������������������       ���Q���?�            �v@"      -                   �?��M���?p           |�@#      *                   �?;��w�?�           �@$      '                   �?�g��m��?�           8�@%      &                   �?��d��?^            �`@������������������������       �      �?Z             `@������������������������       �                     @(      )                   �? 
,�?y           �@������������������������       �@�����?u            `h@������������������������       ��t��G�?           �y@+      ,                   �?��t�k��?"           �}@������������������������       � �ׁsF�?�            �r@������������������������       �u��Q��?q            `f@.      1                   �?���e�?w           Ȃ@/      0                   �?D��ު��?d             f@������������������������       �                     @������������������������       �������?`            �e@������������������������       � �h�7W�?           �z@3      J                   �?�XԐ��?S           �@4      ?                    �?�r����?           0�@5      <                   �?���H��?           �|@6      9                   �?,�+�C�?�            x@7      8                   �?�q�q�?             H@������������������������       ��q�q�?             E@������������������������       �                     @:      ;                   �?X���b�?�            u@������������������������       �        :            �Z@������������������������       ����D�?�            �l@=      >                   �?��c�%�?*            @S@������������������������       �                     @������������������������       �<ݚ)�?'             R@@      G                   �?<�s�F�?�            �y@A      D                   �?�i-x|e�?�            �u@B      C                   �?�q�q�?             E@������������������������       �j���� �?             A@������������������������       �                      @E      F                   �?���}@��?�            �r@������������������������       �`�q�0ܴ?8            �W@������������������������       �,�T�6�?~             j@H      I                   �?     ��?'             P@������������������������       �                     @������������������������       �d��0u��?$             N@K      P                    �?���^���?Q           ��@L      M                   �?��3��?�            `p@������������������������       �                    �K@N      O                   �?.�[%s�?�            �i@������������������������       �D�n�3�?            �L@������������������������       ��7�QJW�?g            �b@Q      R                   �?�:E���?�            `q@������������������������       ����7�?)            �P@S      T                   �?�iʫ{�?�            �j@������������������������       ����3�E�?             J@������������������������       �p=
ף0�?f             d@V      s                   �?�ϐ=p~�?�           X�@W      j                   �?�	��)��?�           ��@X      c                   �?�C����?p           ��@Y      `                   �?�D$}c��?V            @b@Z      ]                    �?X�Հ�+�?N            �`@[      \                   �?��p\�?            �D@������������������������       �                     $@������������������������       ���a�n`�?             ?@^      _                   �?`�q�0ܴ?5            �W@������������������������       � ��WV�?             :@������������������������       � =[y��?%             Q@a      b                    �?���!pc�?             &@������������������������       �և���X�?             @������������������������       �                     @d      g                    �?X�V��[�?           �|@e      f                   �?P�	Q��?y            �h@������������������������       �                     B@������������������������       ���w#'�?`            `d@h      i                   �?8L�0�h�?�            0p@������������������������       � 	��p�?%             M@������������������������       ������?|             i@k      l                   �?h#�.��?9           ��@������������������������       �                    �E@m      p                   �?T$�#���?!           `~@n      o                    �? �|k쭚?�            �r@������������������������       ���:�-�??            @Y@������������������������       ������?u            @i@q      r                    �?D\���;�?m            �f@������������������������       �L�w�=�?-            �Q@������������������������       ��"�*f�?@            @\@t      y                   �?(վH��?#           H�@u      v                   �?h�g%���?g            �e@������������������������       �                     <@w      x                    �?������?Y             b@������������������������       �H�V�e��?&             Q@������������������������       ���c�%�?3            @S@z      {                   �?���?�           ��@������������������������       �                     @|      }                    �?���A�'�?�           ��@������������������������       �vt����?�            Pq@������������������������       ��ת2�%�?           z@      �                   �?�F�*R�?          ���@�      �                    �?v9'�*�?�           Y�@�      �                   �?X؏%���?�           ��@�      �                   �?Z��W(�?
           ��@�      �                   �?|�%�9��?�             y@�      �                   �?���R��?�            �q@�      �                   �?p�)_�5�?�            �m@������������������������       ����^T�?�            `k@������������������������       �@�0�!��?	             1@�      �                   �?
;&����?             G@������������������������       ��n_Y�K�?            �C@������������������������       �                     @�      �                   �? �q�q�?E             ^@������������������������       ����<_�?D            �]@������������������������       �                      @�      �                   �?����?           ��@�      �                   �?��$���?�            �l@�      �                   �? S5W�?t             g@������������������������       � 
�V�?T            �`@������������������������       �                     �I@������������������������       ���<b�ƥ?             G@�      �                   �?�p��K�?�           ��@������������������������       ��e��[�?�            �r@�      �                   �?�.
�XX�?�            �t@������������������������       ��:�^���?X            �`@������������������������       �8EGr��?{             i@�      �                   �?�Ѕ1g��?�           ��@�      �                   �? ܳ�Z�\?�           đ@������������������������       �        �           ��@������������������������       � ��Wnq?0           P}@�      �                   �?�8�ͻ��?�            @w@�      �                   �?��<b���?�            �l@������������������������       ����J�?n            `g@������������������������       �&^�)b�?            �E@������������������������       �.Yd�v��?X            �a@�      �                   �?�pO�?           ��@�      �                   �?�\I7+��?�           �@�      �                   �?j�*�'�?�           �@�      �                   �?����P��?�           Ј@�      �                   �?�1�`jg�?>           �~@������������������������       �h7�z�?*            }@������������������������       ���� ��?             ?@������������������������       ��!5�xi�?�            �r@�      �                   �?Xc!J�ƴ?�            �m@������������������������       �0 �����?V            @^@�      �                   �?�]���?G            �\@������������������������       ��Ń��̧?             E@������������������������       � �й���?+            @R@�      �                   �?����xł?T           ��@�      �                   �?@֊��v�?�           4�@������������������������       � t�)Ї?�           �@������������������������       ����pA�?V            `a@������������������������       �� �Ux?o           x�@�      �                   �?�{Y�'U�?(           �@�      �                   �?���u��?�            �@�      �                   �?N����?�            �u@������������������������       �                     @������������������������       �h!�'nf�?�            0u@�      �                   �?���q��?�            �x@�      �                   �?$V�Ap�?_            �a@������������������������       ��z�G��?             $@������������������������       �pJQg���?X            �`@�      �                   �?�
n�X��?�            `o@������������������������       �r�q��?             @������������������������       �Hm_!'1�?�            �n@�      �                   �?��ؖ��?P           ��@�      �                   �?7�A�0�?�             v@������������������������       �ڡR����?�            `r@������������������������       �l��[B��?$             M@������������������������       ��|R���?s            �g@�      �                   �?h第�?A           (�@�      �                   �?����X��?�            �@�      �                   �?�&/�E�?P             _@�      �                   �?p��@���?3            @U@�      �                    �?Х-��ٹ?+            �R@������������������������       �ܷ��?��?             =@������������������������       ���<b�ƥ?             G@�      �                    �?z�G�z�?             $@������������������������       �                     @������������������������       �      �?             @�      �                    �? ���J��?            �C@������������������������       �        
             (@������������������������       � 7���B�?             ;@�      �                    �?(����?^            �@�      �                   �?�>4ևF�?�             l@������������������������       �V���#�?H            �W@�      �                   �?&X�IN�?Q             `@������������������������       ���V�I��?            �G@������������������������       �v�2t5�?9            �T@�      �                   �?f�Je\��?�            @t@������������������������       ����Y�?e            `d@�      �                   �?֧���?`             d@������������������������       �N1���?#            �N@������������������������       ����ׁs�?=             Y@�      �                   �?@i@��T�?�           ��@�      �                    �?#gI��?           \�@������������������������       ���8Iz»?�           ��@������������������������       ���r����?           ��@�      �                   �?�h.g�;�?�           ��@�      �                    �?H��uӳ?c           Ё@������������������������       �h�����?�             l@������������������������       ���;�?�            �u@�      �                    �?xt~Y�l�?$           @�@������������������������       ���XT梵?�           �@������������������������       ��gߒm��??           |�@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�Bp       h�@     ��@    �W�@     }�@     �@     ��@     P�@     �|@     pz@     `r@     �n@     �i@      f@     �U@     �e@     �U@       @             �X@     �d@      X@     �d@      @             �@     ��@    �6�@     @�@     l�@     ``@     X�@      O@     @�@      F@     �@      F@     �@      @@      _@      �?     �[@      �?      ,@             0�@      ?@     @~@      7@      p@       @      @@      (@              �?      @@      &@     �Q@              @      2@      @      0@       @      (@      �?      @               @      y@     @Q@      ;@      @      7@      @      5@      @       @              @      �?     Pw@      P@      w@      H@     �u@      D@     �t@      D@     �k@      B@     @[@      @      4@              3@       @      0@       @      @              @      0@      @      *@      @      $@      �?      @              @     ��@     P~@     4�@     �q@     ��@     @c@     �X@             Ԥ@     @c@     ��@     @Q@     ��@      "@     <�@      N@     �m@     @U@     Ш@     �_@     �G@             r�@     �_@     Ȧ@      A@     �@      8@     L�@             �@      8@     �}@      $@      f@             pr@      $@     �j@     @W@      d@     �T@     �J@      &@     ��@     �i@     r�@     �U@      �@      @     �@@             ��@      @     H�@      @     0�@      @     �~@      �?     @U@      �?     ė@     @T@      $@             ��@     @T@     P�@     �G@     �@      A@     X�@      :@     @f@       @     Pr@     @]@     �d@      F@      �?             `d@      F@      `@     @R@     @W@      K@      B@      3@     f�@     �@     �r@     �j@     `h@     �Z@     �g@     @T@      f@     @S@      e@     �J@     �W@      A@     �R@      3@       @      8@      *@      @      &@      @      @       @      @       @       @              @      9@              (@      @      *@      @      @               @     �Y@     @[@     @V@      T@     @V@     �N@      T@     �L@     �K@     �H@      9@       @      "@      @      @       @      @       @              3@      *@      =@      *@      7@      @      7@      @                      @     �@     `~@     ��@     `e@     ��@      W@     ��@      @     Pt@      @     0w@      �?      r@             �T@      �?     x�@     �U@     @{@      G@     ؁@     �D@     �y@      ;@      d@      ,@     ��@     �S@     X�@      K@     �p@      @     �q@      I@     �@      9@     �e@      �?      ^@             �K@      �?     �t@      8@     @m@      2@     @X@      @     �{@     �s@      v@     �p@     �k@      c@     ``@      U@     @V@     @Q@     �`@     @\@     �U@     �S@      H@     �A@      W@     �H@      G@      :@      G@      7@     (�@     ��@     �s@     �@     @c@     \�@     �V@     �@      M@      k@              �?      M@     �j@      @      ]@     �I@     �X@     �@@     Px@     �O@     Ѕ@      D@     �j@      @     @b@     �A@     @Q@      7@     0~@      d@     ��@     @X@     �|@              "@     @X@     P|@      @      W@      W@     �v@      H@      R@      F@     r@      P@     ��@       @     �e@      O@      @      @@     �Q@      >@     �z@     �t@     �@     �h@     �@     �\@     H�@      N@     Pw@      @@     @]@             �A@      @@     �T@      <@      p@      K@     �n@      @@     �R@               @      @@      R@       @      D@      >@      @@      6@     @e@      U@     ��@      �?     �V@      �?     �E@             �G@     �T@     ȁ@     �B@     �Z@      :@     �K@      &@     �I@      G@     �|@      6@     �n@      8@     @k@     �`@     <�@     @Q@     �s@     �B@      c@      2@     �K@      @      ;@      *@      <@      3@     @X@      �?     �N@      2@      B@      @@     �d@      @     @Y@       @     �D@      �?      N@      =@     �O@      $@      :@      3@     �B@     �O@     ��@     �D@     �s@      4@     @^@      5@     �h@      6@     Py@      "@      `@               @      "@     �_@      *@     Pq@     �@    ���@     ��@     |�@     ��@     �@      8@     �h@      8@      h@      1@     �F@      1@      3@       @      3@      @      2@      �?      �?      "@                      :@      @     �b@      @     �T@      @     @T@      @     @T@      @              �?      �?              �?      �?                     �P@              @     ��@     ��@     �@     (�@     ��@     ��@     ��@     pt@     `�@     @Q@     �R@      F@      M@      F@      0@             �@      9@      f@      @     y@      4@      I@      p@             �f@      I@     �R@      ]@     �v@     @R@      E@       @      @     �Q@      B@     �E@     0t@     H�@     ��@     ��@     ��@     ��@     @]@     �J@      T@      H@      T@      @             �@     �B@     @h@      �?     �w@      B@      P@     �y@      @     �r@     �N@     �]@     �b@      |@     �_@      I@              @     �_@     �F@      8@      y@     X�@     ��@     ��@      ]@     py@     �K@     Pv@      <@      A@      ,@      <@      ,@      @             0t@      ,@     �Z@              k@      ,@      I@      ;@              @      I@      6@     �u@     �N@     Ps@     �A@      <@      ,@      4@      ,@       @             �q@      5@     �V@      @     �g@      1@      C@      :@              @      C@      6@     @V@     0|@      I@     �j@             �K@      I@     �c@      8@     �@@      :@      _@     �C@     �m@      @     �O@      B@      f@      .@     �B@      5@     `a@     ��@     ܔ@     ��@     �@     `|@     �b@      .@     ``@      @      `@      @      C@              $@      @      <@      @     �V@      �?      9@      @     @P@       @      @      @      @      @             p{@      3@      h@      @      B@             �c@      @     �n@      *@      K@      @      h@      "@     �R@     p|@             �E@     �R@     �y@      @     �r@       @     �X@       @      i@     �Q@     @\@      7@     �G@     �G@     �P@     �a@     І@      Z@     @Q@              <@      Z@     �D@      K@      ,@      I@      ;@     �C@     ��@              @     �C@     x�@      5@      p@      2@     �x@     �@    ���@     >�@     :�@     ��@     x�@     ��@     �y@      M@     �u@     �J@     �l@      ?@     �i@      1@     @i@      ,@      @      6@      8@      .@      8@      @              @     �\@      @     �\@       @             Ȉ@     @Q@     �l@       @      g@      �?     �`@      �?     �I@             �F@      �?     ��@     �P@     pp@     �@@     �r@      A@     �^@      (@     @f@      6@      Y@     �@      �?     ��@             ��@      �?     @}@     �X@     q@      I@     �f@      E@      b@       @     �A@     �H@     @W@     ��@     8�@     �p@     �@     @p@     �@      A@     ��@      ;@     @}@      7@     �{@      @      ;@      @     @r@     @l@      $@     @\@       @     @\@       @     �D@      �?      R@      �?      $@     �@      @     �@      @     ��@      �?     @a@      @     `�@     Њ@     �z@      �@      X@     �q@     �M@      @             �q@     �M@     Pv@     �B@     �_@      0@      @      @      ^@      *@     �l@      5@      @      �?      l@      4@     �j@     �t@     �b@     �i@      ^@     �e@      <@      >@     �P@      _@     ��@     Ӳ@     0u@     �t@      @     @]@      @     �S@      @     �Q@      @      :@      �?     �F@       @       @              @       @       @      �?      C@              (@      �?      :@     �t@      k@     @a@     �U@      P@      ?@     �R@     �K@      :@      5@      H@      A@     @h@     @`@      Y@     �O@     �W@     �P@     �@@      <@     �N@     �C@      p@     ��@     �_@     ��@     �G@     �@     �S@     ��@     �`@     ��@      7@     �@       @      k@      .@     �t@     @[@     ̞@      A@     ��@     �R@     P�@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�B(m         ^                   �?�@�˱��?f           �@       �                    �?2�p|��?�E          @i�@       n                    �?¥"���?�(          @�@                           �?p
E���?�           t�@       
                    �?D^��#��?v           ��@       	                     �?0ζ�_��?t           ��@                            �?�C����?�           x�@������������������������       ��AMĹ�?!            {@������������������������       �"�����?�            �q@������������������������       �r(�܈�?�            pp@������������������������       �                      @       ;                     �? ��:j��?q           ��@       .                    �?�mj����?           a�@                           �?P�HtǪ?�           ��@                           �? G�H- �?�            �p@                           �?���f~%�?�            Pp@                           �?�K}��?�            �i@                           �?�d���?=            �U@������������������������       � qP��B�?<            �U@������������������������       �                     �?������������������������       �        C            @]@������������������������       �        (            �L@                           �?      �?              @������������������������       �                      @������������������������       �                     @       %                    �? #��yA�?H           ��@                            �? ������?B	           ^�@                           �?8��m�>�?M           h�@                           �? ���v��?/           ؋@������������������������       ��~�u��?m           8�@������������������������       �h�kY���?�            @s@������������������������       �H%u��?             I@!       "                    �? �(h�gq?�           �@������������������������       � y����}?u           T�@#       $                    �? :*T�V?�           ��@������������������������       �                   ��@������������������������       � �m�+�?y            @h@&       )                    �?`K]��w�?           ��@'       (                    �?0G���ջ?%             J@������������������������       �z�G�z�?             .@������������������������       �                    �B@*       -                    �?Xa�uYX�?�           T�@+       ,                    �?�;C�ݳ?4           R�@������������������������       � v�/u��?�           h�@������������������������       ��Y B1F�?W           <�@������������������������       ��请���?�            p@/       0                    �?�f� ���?&           p|@������������������������       �                      @1       6                    �?.�*���?$           P|@2       5                    �?���oY��?u            `f@3       4                    �?˒�#�?a            �b@������������������������       �      �?J             \@������������������������       �                     B@������������������������       �¦	^_�?             ?@7       :                    �?���l���?�             q@8       9                    �?@��,*�?�            �m@������������������������       �$�7�L��?X            �a@������������������������       �B�~R(��??            @X@������������������������       �*O���?             B@<       a                    �?p���`��?U	           ^�@=       N                    �?�AJiQ"�?A           &�@>       K                    �?���wMW�?           �z@?       F                    �? +OmT�?�            �x@@       C                    �?�ӭ�a��?�             r@A       B                    �?�E��ӭ�?             B@������������������������       �����X�?            �A@������������������������       �                     �?D       E                    �?�ŇG+��?�            �o@������������������������       �؇���X�?�            �l@������������������������       ����N8�?             5@G       J                    �?PԱ�l�?L            �Z@H       I                    �?`Ӹ����?@            �V@������������������������       �                     @������������������������       �`��F:u�?=            �U@������������������������       �                     1@L       M                    �?�g�y��?             ?@������������������������       ��n_Y�K�?             :@������������������������       �                     @O       ^                    �?�,&A�?/           Ҧ@P       W                    �? �k/�?p           R�@Q       T                    �?� '1�?�           L�@R       S                    �?�++�Qb�?�           �@������������������������       �                     5@������������������������       �@<�Go\�?�           @�@U       V                    �?�4ӏEIp?@           `@������������������������       �                     <@������������������������       � _�	?q?4           �}@X       [                    �?pi����?�           X�@Y       Z                    �?x�+I��?�           ��@������������������������       �                     @������������������������       ��Ռ��?�           ��@\       ]                    �?x�IG�¼?�           ��@������������������������       �                     @������������������������       � "��u�?�           ��@_       `                    �?�z�G��?�             t@������������������������       ��]��?;            �Y@������������������������       �(��6�ռ?�             k@b       c                    �?J��l��?           �y@������������������������       �                     "@d       i                    �?��9jr�?           0y@e       h                    �?��:x�ٳ?�            �h@f       g                    �?4/Gjϵ?c            �c@������������������������       �`����x�?H            �\@������������������������       � �#�Ѵ�?            �E@������������������������       ���Y��]�?            �D@j       m                    �?+`M���?�            �i@k       l                    �?�k���)�?s            �d@������������������������       �d��4�o�?F            �W@������������������������       �r�q��?-             R@������������������������       �p9W��S�?             C@o       �                    �?��ER7w�?�
           U�@p       q                    �?�"A,8�?/           ��@������������������������       ��q�q�?             @r       �                     �?4\�o8�?-           ��@s       ~                    �?6o��޻�?�           L�@t       {                    �?;��i��?6           X�@u       x                    �?`Jj��?�           (�@v       w                    �?x��Q��?�            �l@������������������������       ���^Z��?V            �b@������������������������       �̘SJl��?+            �S@y       z                    �?�ϣ1���?u            �@������������������������       �`���i��?�             v@������������������������       �     ��?�             p@|       }                    �?H�V�e��?@            �Y@������������������������       �h+�v:�?             A@������������������������       �        +             Q@       �                    �?`׀�:M�?�            �r@�       �                    �?���1��?�            �j@������������������������       ���V��;�?l            �d@������������������������       �                    �G@������������������������       ���Y��]�?6            �T@�       �                    �?���:VW�?6           P�@�       �                    �?��*���?�           ��@�       �                    �?o׭��?b            �b@�       �                    �?�Cc}h,�?J             \@������������������������       �LMc����?6            @T@������������������������       ��4�����?             ?@������������������������       ����@��?            �B@�       �                    �?0���|�?$            |@�       �                    �? Ud2h�?           @y@������������������������       �@��O�A�?�            �q@������������������������       �P����?T            �]@������������������������       ����.�6�?             G@�       �                    �?`��4Eѓ?�            0s@�       �                    �?�6H�Z�?�            @m@������������������������       ��q�q�?l             h@������������������������       �                     E@������������������������       � �й���?+            @R@�       �                    �?~��+߆�?�           �@�       �                    �?� �a��?�           H�@�       �                     �?h�3S<��?           �@�       �                    �?���8�5�?0           }@������������������������       �      �?              @������������������������       �H�����?+           �|@�       �                    �?4Qi0���?�            w@������������������������       �                     @������������������������       ��C��2(�?�            �v@�       �                     �?�B�����?�             j@������������������������       �z8,���?V             _@������������������������       ��P�����?5             U@�       �                    �?lQ���?!           ��@�       �                    �?�҉9��?           `�@�       �                     �?���J�?�           0�@�       �                    �?��ҘR�?            {@������������������������       ��q�q�?             @������������������������       �DI�o��?           �z@�       �                    �?�c:��?�            @q@������������������������       �8�Z$���?             *@������������������������       �p-*<�(�?�            pp@�       �                     �?P�~D&�?S            �`@������������������������       �l�Ӑ���?6            �U@������������������������       �t/*�?            �G@�       �                    �?�P#��6�?           py@�       �                     �?8���u�?�            `s@�       �                    �?L�'��T�?{            @f@������������������������       �                     @������������������������       �p}"����?y            �e@�       �                    �?���7�?R            �`@������������������������       �                      @������������������������       �Hn�.P��?N             _@�       �                     �?�E���?>            @X@������������������������       ����b���?#            �L@������������������������       ��G�z�?             D@�                          �?�����?�           ��@�       �                    �?4��N�0�?�
           +�@�       �                    �?�-��Y�?            ��@�       �                    �?F�-��?s           6�@�       �                    �?ڡR����?           �{@�       �                    �?��W3�?�            0v@�       �                     �?     \�?K             `@������������������������       �8�A�0��?             6@������������������������       ��&=�w��?;            �Z@�       �                     �?�t�����?�            `l@�       �                    �?(Q����?D            @Y@������������������������       �,�|%�v�?7            @U@������������������������       �                     0@�       �                    �?�ՙ/�?U            �_@������������������������       �Z��Yo��?S             _@������������������������       �                      @�       �                    �?�a7���?:            �U@�       �                     �?�,�٧��?3            �S@�       �                    �?:	��ʵ�?            �F@������������������������       ��q�q�?             @������������������������       �r�q��?             E@�       �                    �?�!���?             A@������������������������       �                     @������������������������       �d��0u��?             >@������������������������       �                     @�       �                    �? ��9K�?U           ��@�       �                    �?�T
�8�?Y           x�@�       �                     �?�4�j�ǡ?�            �x@�       �                    �?�S\��?             k@������������������������       �                      @������������������������       ��ɻ9�?z             j@�       �                    �?�Y�ߠ?v            `f@������������������������       �                      @������������������������       �P����?u             f@�       �                    �?�dJ�Ҙ?d            `d@������������������������       �                     @�       �                     �?�Fǌ��?a            �c@������������������������       �        6             W@������������������������       �Pa�	�?+            �P@�       �                    �?�u�%j�?�           ̒@�       �                    �?������?�           ��@������������������������       �                      @�       �                     �?����̺?�           Ј@������������������������       ��*v��?�            @x@������������������������       �������?�            `y@�       �                     �?̐� �?           py@������������������������       �`.��A��?�            �m@������������������������       �4և����?l             e@�       �                    �?��
��?�           �@�       �                    �? ��7h)�?�           ��@�       �                    �? [ ɪ�?e           ��@������������������������       �        1            �T@�       �                     �?`ar	��?4           `~@������������������������       ���S����?z            �g@������������������������       ���F�D�?�            �r@�       �                     �?�K}��?D            �Y@�       �                    �?P�Lt�<�?             C@������������������������       �                      @������������������������       �������?             B@������������������������       �        (             P@�       �                    �?n� ��?           Pz@�       �                     �?��רi�?�            �s@������������������������       �6DSbq��?P             a@������������������������       �:���W�?v             f@�       �                     �?�m��Wv�?>             [@������������������������       ��BE����?"             O@������������������������       �\X��t�?             G@�       
                    �?@,�.���?�           4�@�                          �?V�����?&           �|@�                          �?Rq�����?�            �o@�       �                    �?t���D�?8            �U@������������������������       �                     @                          �?��Q���?3             T@������������������������       ���� ��?             ?@������������������������       �                    �H@                         �? 
��р�?n             e@������������������������       �r�q��?             @������������������������       �8$�s���?j            `d@                         �?D|U��@�?�             i@������������������������       �                     "@      	                   �?     ��?y             h@������������������������       �������?E             [@������������������������       ���X��?4             U@                         �?�S�V@��?�           (�@                         �?N�W+U�?�            v@                         �?�q�q�?S             ^@                         �? >�֕�?4            �Q@������������������������       ��IєX�?             1@������������������������       � �h�7W�?%            �J@������������������������       �HP�s��?             I@                         �?@|����?�             m@������������������������       �                     ?@������������������������       ��M����?}            @i@                         �?�48X'�?�            @r@                         �?���"F��?�            `i@������������������������       �                     @������������������������       � �M*k�?�            �h@������������������������       ���=���?;            @V@      ;                   �?̄/���?�           =�@      2                   �? ��=���?l           ��@      +                   �?|����e�?           ��@      $                    �?��S��?�           �@      !                   �?��o	��?!            }@                          �?6#�����?�            w@������������������������       �8��%���?�            �m@������������������������       �0�!F��?R            �`@"      #                   �?���c��?=            �W@������������������������       ��d�����?             C@������������������������       �        $            �L@%      (                   �?Jo�~�M�?�           ��@&      '                   �?�IєX�?M           x�@������������������������       �xWT�Nt�?9           �~@������������������������       �<���D�?            �@@)      *                   �?�S�A�?g            �d@������������������������       �hx<?v��?L            �]@������������������������       �=QcG��?            �G@,      /                    �?t����?7           0@-      .                   �?�C$���?d             c@������������������������       ��1e�3��?M            �]@������������������������       ���?^�k�?            �A@0      1                   �?�'#"�o�?�            �u@������������������������       ��==Q�P�?�            �q@������������������������       ���v$���?$            �N@3      8                   �?��Mx?`           B�@4      7                   �?����v9v?�           ��@5      6                    �? ��ϰ`y?           $�@������������������������       � yqn�{?~           @�@������������������������       ��7A|
�w?�           �@������������������������       �        �            �l@9      :                    �?�� �U�z?�           ̗@������������������������       ����H��?            �}@������������������������       � ��]�xw?�           P�@<      G                   �?n���?�           H�@=      B                    �?�����g�?�           ��@>      A                   �?���i@�?'           �{@?      @                   �?�
0����?�            �q@������������������������       �r�q��?             @������������������������       ���27
��?�            `q@������������������������       ���絹�?o            `d@C      F                   �?�[���?w           ��@D      E                   �?$M���?�            `t@������������������������       ����Q��?             $@������������������������       ��+ت�M�?�            �s@������������������������       �
���?�            @n@H      W                   �?"�G�6�?�           ��@I      P                   �?|I���?�           ��@J      M                    �?�E�0�/�?�             s@K      L                   �?ཕvt�?a            �b@������������������������       ������H�?             "@������������������������       �hA� �?\            �a@N      O                   �?��a�n`�?_            `c@������������������������       �                     @������������������������       �46��e-�?[            �b@Q      T                    �?H���?           |@R      S                   �?ףp=
�?z            �g@������������������������       �                      @������������������������       � .2��A�?x            �g@U      V                   �?�MI8d�?�            0p@������������������������       ��<ݚ�?             "@������������������������       ��J�4�?�            @o@X      [                    �?����-�?           �{@Y      Z                   �?��+�ޯ�?u            �f@������������������������       ��~8�e�?            �I@������������������������       ���^@=��?X            ``@\      ]                   �?~4y�_R�?�            `p@������������������������       ���WV��?#             J@������������������������       �<=�,S��?w            @j@_      �                   �? >1M��?W           ���@`      �                   �?j"e��?Y           X�@a      r                    �?z��bss�?G           ��@b      m                   �?`�Cb؟�?�           ��@c      h                   �?^
`,���?�           ��@d      g                   �?@��MP��?�           ��@e      f                   �?ė����?�            ps@������������������������       �ףp=
�?             $@������������������������       �^����?�            �r@������������������������       ��䖑��?�            �w@i      l                   �?(�>m�C�?8            @j      k                   �?(֌��)�?�            `p@������������������������       ����Q��?             @������������������������       ��U�'���?�            p@������������������������       �8��%���?�            �m@n      q                   �?�4F����?�            �i@o      p                   �?8^s]e�?&             M@������������������������       �      �?              @������������������������       ��-���?"             I@������������������������       ���m.	�?d            `b@s      �                   �?��j�9�?�           h�@t      }                   �?�E'�>�?@           ��@u      z                   �?�v�M��?Y           H�@v      w                   �?P��MO�?�             o@������������������������       �                     @x      y                   �?`[�͏�?�            �n@������������������������       ����y4F�?	             3@������������������������       �D��_$�?�            @l@{      |                   �?R��Xp�?�             s@������������������������       �                     �?������������������������       �:@�r{�?�            �r@~      �                   �?���]P0�?�            �v@      �                   �?zv�X��?o             f@������������������������       �                      @������������������������       �T����1�?m            �e@������������������������       �@-�_ .�?x             g@�      �                   �?|�Pk��?~             i@������������������������       �                      @�      �                   �?J������?}            �h@�      �                   �?�	j*D�?#             J@������������������������       �                      @������������������������       � �o_��?!             I@������������������������       ��c!�^�?Z            @b@�      �                   �?"�ܕ���?           �@������������������������       �        
             2@�      �                    �?.\r����?           ��@�      �                   �?���+�?�           ��@�      �                   �?_U/2�?�            �p@�      �                   �?���N8�?             5@������������������������       �ףp=
�?             $@������������������������       �                     &@�      �                   �?$H�fpM�?�            �n@�      �                   �?�Ha�3�?|            `h@������������������������       �2�[���?R            �_@������������������������       ��t����?*             Q@������������������������       � s�n_Y�?"             J@�      �                   �?L�'�7��?           ��@�      �                   �?���zS��?P           ��@������������������������       ��7���?�            @w@������������������������       �(32v�c�?`            `d@������������������������       �h>#j�x�?�            �q@�      �                   �?���n��?X           ��@�      �                   �?Z'8of�?           �@�      �                   �?T)�b�w�?�             l@�      �                   �?�����H�?             2@������������������������       �8�Z$���?             *@������������������������       �                     @�      �                   �?������?�            �i@������������������������       ��L�w��?Y            �a@������������������������       ����`��?+            �P@�      �                   �?�Ber�J�?}           �@������������������������       ��Y\��޽?            {@������������������������       �T���D9�?n            �e@�      �                   �?p��tKn�?L           �@�      �                   �?�):u��?6            @S@������������������������       �                      @������������������������       ���x�5��?0            @Q@������������������������       �He��+��?           �z@�      �                   �?��"����?�           �@�      �                   �?>��wff�?l           ֳ@�      �                   �?�媀]�?�           ��@�      �                   �?f���?           �@�      �                    �?.T�߸��?�            @w@�      �                   �?�������?�             h@������������������������       �                     &@������������������������       ��-�c��?x            �f@�      �                   �?�/��(�?k            `f@������������������������       �                     &@������������������������       ��ՙ/�?d             e@�      �                    �?x�ǋ��?3           ��@������������������������       �XP���Ƿ?&           p}@������������������������       ����g�X�?           �{@�      �                    �?��xy�?�           ��@�      �                   �?P�X���?Y           ��@�      �                   �?������?S             `@������������������������       �"pc�
�?             6@������������������������       �ʫe�s,�?E            �Z@������������������������       ��x�?���?           ؉@�      �                   �?æ�!F�?r           4�@�      �                   �?�G��l��?�            @j@������������������������       � ���J��?            �C@������������������������       �D�n�3�?g            `e@������������������������       �PU��?�           �@�      �                   �?�aV����?�           $�@�      �                   �?���D�?�           ��@�      �                    �?�/jF�[�?�            �n@�      �                   �?���A��?e            �b@������������������������       �                     @������������������������       ���ӭ�a�?b             b@�      �                   �?v�C��?=            �X@������������������������       �                     $@������������������������       �:��?7            @V@�      �                    �?H�\Qg	�?)           �}@������������������������       �����a�?�            �n@������������������������       �3e��?�            `m@�      �                   �?@s�RF�?�           ��@�      �                   �?@lܯ ��?J            �]@�      �                    �?      �?             0@������������������������       �                     $@������������������������       ��q�q�?             @�      �                    �?��>��?B            �Y@������������������������       ��lg����?            �E@������������������������       �*;L]n�?'             N@�      �                    �?���7�?n           ��@������������������������       ���s�n�?�             j@������������������������       ��ȉo(��?�            �v@�      �                   �?�
�b���?�           *�@�      �                   �?Ċ����?           �z@�      �                    �?D]��;��?s            @h@�      �                   �?��a����?4            �T@������������������������       �                     �?������������������������       ��p ��?3            �T@�      �                   �?|$�����??            �[@������������������������       �                     0@������������������������       ��\��N��?7            �W@�      �                    �? ��X��?�            �m@�      �                   �?���
��?>            �Z@������������������������       �ףp=
�?             4@������������������������       ��(~�[�?3            �U@�      �                   �?B@��S��?V             `@������������������������       ��IєX�?             A@������������������������       ��\��N��?>            �W@�      �                   �?��9 h۵?�           Τ@�      �                    �?X#o2�?A           ��@������������������������       �XY��p9�?�             n@������������������������       ��Iч�r�?�            r@�      �                    �?M#�w@�?J           ��@������������������������       ���gU?n�?�           ��@������������������������       �P>CZ���?^           �@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B0       ^�@     ��@    ���@     �@    ���@     $�@     ��@     H�@     ��@     �|@     p�@     �|@     �z@      r@     �m@     �h@     `h@      W@     �W@      e@       @             ��@     (�@     @�@     �@     �@     �f@     �p@      @     0p@       @     @i@       @     @U@       @      U@       @      �?             @]@             �L@              @       @               @      @             ڸ@     `f@     �@     �L@     Ћ@     �I@     p�@     �F@     8�@      @@     pr@      *@      F@      @     ��@      @     @�@      @     ��@      �?     ��@              h@      �?     Ȥ@     �^@     �H@      @      (@      @     �B@             f�@     �]@     ��@      Y@     ��@      J@     |�@      H@     �m@      3@     @W@     �v@               @     @W@     �v@      0@     `d@      @     �a@      @     @Z@              B@      "@      6@     @S@     �h@      P@     �e@     �B@      Z@      ;@     �Q@      *@      7@     ��@     �~@     ڨ@     �d@     �v@      P@     �u@      H@     �n@      F@      :@      $@      9@      $@      �?             @k@      A@     �h@     �@@      4@      �?     �Y@      @     �U@      @      @             �T@      @      1@              .@      0@      $@      0@      @             �@     �Y@     ��@     @U@     4�@      @     ��@      @      5@             �@      @     P@      �?      <@             �}@      �?     �@     �S@     ��@     �B@      @             h�@     �B@     ��@      E@      @             ��@      E@     �r@      1@     �X@      @     �i@      *@     @V@     0t@              "@     @V@     �s@       @     �g@      @     �b@      @     @[@       @     �D@      �?      D@     @T@      _@     �Q@     @X@     �B@      M@     �@@     �C@      &@      ;@     *�@      �@     ��@     ��@       @      �?     ��@     ��@      �@     �v@      �@     �R@     x�@      K@      g@      F@     @^@      =@      P@      .@     ��@      $@     �u@       @     �o@       @     @T@      5@      *@      5@      Q@              @     @r@       @     �j@       @     �d@             �G@       @      T@     0�@     @x@     �@      U@     @R@      S@     @P@     �G@      F@     �B@      5@      $@       @      =@     �{@       @     �x@      @     �q@      @      ]@       @     �E@      @      @      s@       @      m@       @     �g@              E@      �?      R@     ��@     �|@     ȉ@      k@     ؇@     �Q@     �z@      C@      @      @     pz@      A@      u@     �@@      @             �t@     �@@      O@     @b@     �B@     �U@      9@     �M@     ��@     `n@     H�@     `d@     (�@     @P@     `x@      F@       @      �?     @x@     �E@     �o@      5@      &@       @     �n@      3@      B@     �X@      <@     �M@       @     �C@     pt@      T@     0r@      3@     �d@      *@      @             @d@      *@     �_@      @       @             �]@      @      B@     �N@      7@      A@      *@      ;@     �@     ��@     �@     ��@     ��@     �@     ��@     �u@     �f@     Pp@     @_@     �l@      *@     �\@      "@      *@      @     �Y@      \@     �\@      P@     �B@      H@     �B@      0@              H@     �S@      G@     �S@       @             �K@      ?@      H@      ?@     �B@       @       @      �?     �A@      @      &@      7@              @      &@      3@      @             (�@      V@     0�@      "@     Px@      @     �j@      @       @             �i@      @      f@      @       @             �e@      @      d@       @      @             �c@       @      W@              P@       @     ��@     �S@     ��@      F@       @             p�@      F@     �v@      8@      x@      4@     @w@     �A@     `k@      4@      c@      .@     �d@     ��@       @     ��@      @     ��@             �T@      @     �}@      �?     �g@      @     0r@      �?     @Y@      �?     �B@               @      �?     �A@              P@     �c@     `p@      \@      i@     �H@     �U@     �O@     �\@     �G@     �N@      5@     �D@      :@      4@     p�@     ��@     @n@     �j@     �j@     �E@     �J@     �@@              @     �J@      ;@      @      ;@     �H@             �c@      $@      @      �?     @c@      "@      >@     `e@              "@      >@     @d@      @     @Z@      ;@     �L@     �q@     �v@     �J@     �r@      I@     �Q@      @     �P@      �?      0@      @      I@      G@      @      @     �l@              ?@      @     �h@     �l@     �N@     `g@      0@      @             �f@      0@      F@     �F@     ��@     P�@     `�@     ��@     �@     ؑ@     @y@     ��@      k@      o@     �b@     �k@      5@     �j@      `@      @     �P@      <@      $@      <@     �L@             �g@     �@      ?@      @      ;@     0}@      @      =@     �c@      "@     @\@      @      F@      @     �[@     Px@     �D@      \@      @     �[@      A@      �?     @Q@     Pq@      "@     @q@      N@      �?      $@     .�@      @     ��@      @     �@       @     0�@      @     ��@             �l@      @     ��@       @     �}@      @     D�@     ��@     �@     `�@     �v@     r@     �c@     �o@      ?@      @      �?      o@      >@      B@     �_@     �v@     �i@     �q@      F@      @      @     @q@      D@     @T@      d@     ��@     �u@     ��@     �T@     �q@      6@     �a@      @       @      �?     �`@      @     �a@      .@      @             �`@      .@     @x@     �N@     `e@      3@       @              e@      3@      k@      E@      @       @     @j@      D@     �f@     Pp@     �T@      Y@      6@      =@      N@     �Q@     @Y@      d@      7@      =@     �S@     �`@     ڣ@     ��@     Е@     ȫ@     �@     �@     �@     ��@     �{@     H�@     @o@     `{@     @k@     @W@      �?      "@      k@      U@      @@     �u@     �g@     0s@     @e@      W@       @      @      e@     @V@      5@     �j@     @P@     �a@      D@      2@      @      @     �B@      *@      9@     �^@     �x@     ��@     �u@     ��@     �k@     �t@      f@      R@      @             �e@      R@      @      .@      e@     �L@      G@      p@              �?      G@     p@     �_@     @m@     @]@     �M@               @     @]@     �L@      $@     �e@     �E@     �c@               @     �E@     `c@      B@      0@               @      B@      ,@      @     `a@     @     x�@              2@     @     0�@      p@     �@     �f@     �U@      �?      4@      �?      "@              &@     �f@     �P@     `a@      L@     �V@      B@      H@      4@     �D@      &@     @S@     0�@      H@     p~@     �@@     0u@      .@     �b@      =@     �o@     �m@     <�@      f@     ��@     �_@     �X@       @      0@       @      &@              @     @_@     �T@     @V@     �I@      B@      ?@      I@     x�@      ;@     py@      7@      c@      O@     �{@     �D@      B@               @     �D@      <@      5@     �y@     �@     r�@     ��@     ��@     8�@     L�@      o@     0�@      i@     `e@     @X@      X@              &@     @X@     @U@      Z@     �R@              &@      Z@      P@     �G@     �@      7@      |@      8@     z@     �r@     4�@     @a@     ��@      S@     �J@      @      2@      R@     �A@      O@     �@     �d@     ��@      Y@     �[@      �?      C@     �X@      R@     @P@     �@     q@     ��@     �f@      �@     �a@     �Z@     �T@     �P@              @     �T@      O@     �M@      D@              $@     �M@      >@     �D@     `{@      3@      l@      6@     �j@     �V@     ��@     @P@      K@      @      (@              $@      @       @     �N@      E@      ;@      0@      A@      :@      :@     �@      $@     �h@      0@     �u@     t@     ��@     @i@     �l@      W@     �Y@      E@     �D@              �?      E@      D@      I@     �N@              0@      I@     �F@     �[@     �_@      M@     �H@       @      2@      L@      ?@      J@     @S@       @      @@      I@     �F@     �]@     �@      ?@     0@      (@     �l@      3@     �p@      V@     ��@      B@     `�@      J@     D�@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�B(m         �                    �?b�/=��?�e           �@       �                    �?�w����?�5           B�@       T                    �?0ռ[~�?�(          �(�@                           �?��N�j�?r           ��@                           �?􆧽u��?`           ��@                            �?������?_           ��@       
                    �?����?�           ��@       	                     �?�-�Z�?�           ��@������������������������       ���A����?           0z@������������������������       �b;
!��?�            0s@������������������������       �                     �?                           �?6Pc���?�            �k@������������������������       � �a�e��?�            �k@������������������������       �                     �?������������������������       �                      @       =                    �?��[:���?           :�@                           �?�?�(|�?�           ��@                            �?XB���?^             b@                           �?Ц�f*�?H            �[@                           �?����q�?G            @[@������������������������       �����?�?<            �V@������������������������       �                     3@������������������������       �                     �?                           �? >�֕�?            �A@������������������������       �(;L]n�?             >@������������������������       �z�G�z�?             @       ,                     �?�2�`XH�?w           d�@       '                    �?��S�ۿ?j           h�@       $                    �?��}S߷?Z           ��@       !                    �?�e ��5�?8           Ќ@                            �?Ю�-(�?m           ��@������������������������       �8��"s�?\           (�@������������������������       �`2U0*��?             9@"       #                    �?��҂� �?�            �u@������������������������       � �˟?�            �s@������������������������       �                     ?@%       &                    �?���y4F�?"            �L@������������������������       ��T`�[k�?            �J@������������������������       �                     @(       )                    �?R�}e�.�?             :@������������������������       �؇���X�?             ,@*       +                    �?�q�q�?             (@������������������������       �X�<ݚ�?             "@������������������������       ��q�q�?             @-       8                    �?R,RMn�?           �z@.       3                    �?T}_���?�             w@/       2                    �?d�6��:�?�            @o@0       1                    �?��
Bo5�?�            @n@������������������������       �*
;&���?�            �l@������������������������       ��8��8��?             (@������������������������       �      �?              @4       7                    �?�(\����?K             ^@5       6                    �? �w5�?J            �]@������������������������       �`�LVXz�?A            �X@������������������������       �        	             3@������������������������       �                      @9       <                    �?П[;U��?              M@:       ;                    �?Np�����?            �I@������������������������       �X�<ݚ�?            �F@������������������������       �                     @������������������������       �                     @>       S                    �?~���]c�?=           0@?       N                    �?6��z��?!           `|@@       G                    �?�q5�U�?�            `x@A       D                     �?�1���?�            @n@B       C                    �?�����?a            �b@������������������������       ���+7��?[            @a@������������������������       �      �?             $@E       F                    �?z�J��?B            �W@������������������������       ���S���??            �V@������������������������       �                     @H       K                    �?����>�?T            �b@I       J                     �?
��[��?I            @`@������������������������       �NKF����?3            @V@������������������������       �D^��#��?            �D@L       M                     �?�<ݚ�?             2@������������������������       �����X�?             @������������������������       �"pc�
�?             &@O       P                     �?     x�?*             P@������������������������       �؀�:M�?            �B@Q       R                    �?�q�q�?             ;@������������������������       ���<b���?             7@������������������������       �                     @������������������������       �                    �F@U       �                    �? �ی�B�?U!           g�@V       �                    �?��(�p �?�          ���@W       t                    �?�lӋ�?�           ��@X       e                    �?�'��f�?�           /�@Y       `                    �?@�t#�?�	           ��@Z       ]                     �?�vp I��?]           �@[       \                    �?��"���?�           ��@������������������������       �        C             Z@������������������������       � {��Y��?q           @�@^       _                    �? ž��?�           ��@������������������������       �        
             ,@������������������������       � g�yB�?�           (�@a       b                    �? <S�(�Q?`           �@������������������������       �        !             K@c       d                     �? �$�R??           <�@������������������������       �        	           ��@������������������������       ��ȲA��p?6           �~@f       m                     �?������?�	           ��@g       j                    �?�%`)���?]           �@h       i                    �?:-�5��?�           l�@������������������������       �                     @������������������������       �ȫ�0�?�           `�@k       l                    �?�^�� �?i           T�@������������������������       �                     �?������������������������       ��	:6&�?h           P�@n       q                    �?��L��u�?x           ��@o       p                    �?����|��?�            �@������������������������       �                     @������������������������       ��qqa���?�           Ѕ@r       s                    �?�yr�?c�?�           x�@������������������������       �                     @������������������������       ��Y�ɖ�?�           P�@u       |                    �?��F%���?S           �@v       y                    �?@
�J�?�           ��@w       x                     �? f(<��?�           ؂@������������������������       �@�s���?�            �u@������������������������       �`���£?�            �o@z       {                     �?��*X�u?�            �w@������������������������       ��}.yI�?�            �k@������������������������       �        _            `c@}       �                     �?�����?�           p�@~                           �?l���	�?J           �@������������������������       �l��.���?$           0}@������������������������       ���D�܇�?&           �~@�       �                    �?�s�й�?�           ��@������������������������       ��2(&��?�             v@������������������������       �0�|#�p�?�            �o@�       �                    �?`��F:u�?�           ��@�       �                    �? �qǩ�?�            �@�       �                    �? tly47{?�            �r@������������������������       �                     @�       �                     �? 7O�W}{?�            �r@������������������������       �@_�M�q�?k            �g@������������������������       �        C            �Z@�       �                     �?��)�G��?'           @}@������������������������       �     ��?�             p@������������������������       ��NW���?�            �j@�       �                    �?����&!�?�            �v@�       �                     �?@��!�Q�?J            @Z@������������������������       �        (            �N@������������������������       �`���i��?"             F@�       �                     �?֨!t��?�             p@������������������������       ��K�	H�?l             c@������������������������       ���?^�k�??            @Z@�       �                    �?jX?����?�           �@�       �                    �?ʐ��VS�?�           ��@�       �                     �?P-{ R�?`           �@������������������������       ����f+�?�            `u@������������������������       ��L��?�            `i@�       �                    �?D|X\�G�?G           p�@�       �                     �?j�Je���?�            �x@������������������������       �xk�9�?�            `m@������������������������       ��Hvk��?]            �c@�       �                     �?:-�.A�?V            �`@������������������������       �v���EO�?/            �Q@������������������������       ��q�q�?'            �O@�       �                    �?<c��.�?�           ��@�       �                     �?\��Ho�?�           ��@�       �                    �?b�+����?�            �v@������������������������       �<K���m�?�            `g@������������������������       �{�����?k            �e@�       �                    �?k��9�?�            �p@������������������������       �B��c�?e            `e@������������������������       ��"���r�?A            �X@�       �                     �?����3��?j            �c@������������������������       ����|���?2            @S@������������������������       �t�C�#��?8            �S@�       �                    �?h�B�H��?�           e�@�       �                     �?�O�Af<�?�           X�@�       �                    �?�#N|ї�?X           ��@�       �                    �?�Y����?I           �@������������������������       �                     �?�       �                    �?6@����?H           �@�       �                    �?�Ʈ�?           0{@�       �                    �?��3EaǼ?r             g@������������������������       �$�q-�?Z            �a@������������������������       �                    �D@�       �                    �?����T�?�            `o@������������������������       ����=A�?`             c@������������������������       ��q�q�?F            �X@�       �                    �?ޚ)�?0             R@������������������������       �     ��?             @@������������������������       ����Q��?             D@�       �                    �?�5e�U!�?           (�@�       �                    �?P����?�           ��@������������������������       ��u����?           �y@������������������������       ���L�J2�?�            �o@������������������������       �t/*�?a            �a@�       �                    �?��T��?�           ,�@�       �                    �?�\ڋ�?�           ��@�       �                    �?��^��~�?R           ��@�       �                    �?Pns��ޭ?P            �`@������������������������       �                     @������������������������       ��i�y�?K            �_@�       �                    �?"pc�
�?           �x@������������������������       �r�0?��?F            �Z@�       �                    �?�e!p���?�            r@������������������������       �                      @������������������������       �����?�            �q@�       �                    �?     ��?�             p@������������������������       �                     �?�       �                    �?�G�c��?�            �o@�       �                    �?
�c�Z�?A             Y@������������������������       ���Y��]�?            �D@������������������������       ��ݜ����?)            �M@������������������������       ���F��?e            `c@�       �                    �?������?�            @o@������������������������       �                     �?�       �                    �?�}#���?�             o@�       �                    �?�*v��?9            @X@������������������������       � ��WV�?              J@������������������������       ���Hg���?            �F@������������������������       ��}�+r��?S             c@�       �                    �?��C�L��?           r�@�       �                    �?�ů��6�?/           .�@�       �                     �? f��L��?�           $�@�       �                    �?�?����?�           8�@������������������������       �        a            �b@�       �                    �?�a�OR�?�           ��@������������������������       ��q�q�?L            �^@������������������������       ��0�Z��?6           `}@�       �                    �?�Nh��?�           �@������������������������       �`���i��?X            �`@�       �                    �?�s�M�L�?Q           ��@������������������������       ��������?8             V@������������������������       �`�F���?           `|@�       �                     �?̹� &��?�           p�@�       �                    �?dk�����?�             u@�       �                    �?�N�#/�?U            @`@������������������������       �        "             M@������������������������       �P��E��?3             R@������������������������       �b �57�?�            �i@�       �                    �?D���D|�?�            �s@������������������������       �                     E@�       �                    �?<���|��?�            @q@������������������������       �6YE�t�?            �@@������������������������       �������?�            `n@�       �                    �?�N��#��?�           �@�       �                     �?��L�J2�?�            �o@�       �                    �?�?�0�!�?S             a@������������������������       �`��>�ϗ?2            @U@������������������������       �������?!            �I@�       �                    �?�ݜ�?K            @]@������������������������       �P�2E��?)            @P@������������������������       ��θ�?"             J@�       �                     �?xRdΕ�?R           (�@������������������������       ���GEI_�?�            �n@������������������������       ����n4s�?�            s@�       �                   �?`���OP�?60           ��@�       _                   �?�Jq�m�?�           h�@�       >                   �?
����?           �@       /                   �?:,�i��?�           ��@                         �?P��j�?t           8�@                         �?�7娩�?�           ��@                         �?
�r13G�?�            �u@                          �?�8��8N�?7             X@������������������������       ������?             3@������������������������       ��e���@�?*            @S@      
                    �?���t!V�?�            @o@      	                   �?n�tl��??            �Z@������������������������       ���̅��?8            �W@������������������������       �                     (@                         �?zng���?Z            �a@������������������������       �`n��k��?W            `a@������������������������       �                     @                         �?�9�3+�?�           $�@                          �?`8�.��?�             w@                         �? r���?�            �g@������������������������       �                     @������������������������       �@�Gpm��?}             g@                         �? �.�?Ƞ?s            �f@������������������������       �                     �?������������������������       ��Y�ߠ?r            `f@                          �?�E����?�           ��@������������������������       � fM6��?�            px@������������������������       � �lV}�?�             y@      (                   �?�θn��?�           ȅ@      !                    �?     ��?�             p@                         �?,�d�vK�?\            �a@                         �?      �?             @������������������������       �      �?              @������������������������       �                      @                          �?D��*�4�?X            @a@������������������������       �z�G�z�?             I@������������������������       �        =             V@"      %                   �?F�t�K��?N            �\@#      $                   �?���Q��?            �A@������������������������       �                     �?������������������������       �j���� �?             A@&      '                   �?�Fǌ��?5            �S@������������������������       �                     �?������������������������       ��(�Tw�?4            �S@)      ,                    �?�ڇ��*�?           �{@*      +                   �?Xl���?�            �l@������������������������       �                     @������������������������       �      �?�             l@-      .                   �?�J�T�?�            �j@������������������������       �                     @������������������������       ���?^�k�?�            @j@0      7                   �?L񙤁�?           �{@1      4                    �?�g�W��?�            Ps@2      3                   �?F��ӭ��?V             b@������������������������       �`2U0*��?             9@������������������������       ��n\�GZ�?I            �]@5      6                   �?�q�q�?f            �d@������������������������       ��r����?	             .@������������������������       � �o_��?]            �b@8      ;                    �?Pa�.l�?U            �`@9      :                   �?���;+"�?.            �S@������������������������       �                     @������������������������       ���T���?+            @R@<      =                   �?�eP*L��?'            �K@������������������������       �                     @������������������������       �`�(c�?$            �H@?      L                   �?ȵHPS!�?�           x�@@      G                    �?@��v�?�           ��@A      D                   �? �w5�?�            �m@B      C                   �?@_�M�q�?            �g@������������������������       �                     4@������������������������       �@c����?s            @e@E      F                   �?��<b�ƥ?             G@������������������������       �                     @������������������������       � qP��B�?            �E@H      K                   �?�+#߿��?	           �z@I      J                   �?����|��?�             v@������������������������       �        +            �R@������������������������       ��̳n�?�            `q@������������������������       ��?�|�?)            �R@M      T                   �?v]FN��?�           ��@N      Q                    �?6DSbq��?�            �y@O      P                   �?��n�u�?f            �f@������������������������       ��m���?D            �]@������������������������       �b����?"            �O@R      S                   �?|x$���?�            `l@������������������������       �v���?s             f@������������������������       �H.�!���?             I@U      \                   �?HF�{o�?�           8�@V      Y                    �?��j�?            �@W      X                   �?8��8��?            x@������������������������       �                     �?������������������������       ���`�]��?           �w@Z      [                   �?0g�BJ��?           @|@������������������������       �                     @������������������������       �8և����?            |@]      ^                    �?�)x��?�            �t@������������������������       �$��$�L�?g            �c@������������������������       ����tT��?j            �e@`      �                   �?F_G���?�           ��@a      v                   �?�������?<           ��@b      k                    �?�Y����?^           2�@c      j                   �?a" @n�?�           |�@d      g                   �?�d�Ì��?           �x@e      f                   �?���9���?�            �s@������������������������       ����x��?�            �i@������������������������       ��g+��@�?H            �[@h      i                   �?NP�<��?:            �T@������������������������       �$�q-�?             :@������������������������       ����U�?'            �L@������������������������       �        �           ��@l      q                   �?��*�?�           �@m      p                   �?�Vy��?*           h�@n      o                   �?��!���?�           ��@������������������������       �@[p��ж?6           �~@������������������������       ���?^�k�?U            �a@������������������������       � 9���n?�           ��@r      u                   �?�X�#�?�             l@s      t                   �?��ӭ�a�?0             R@������������������������       �r�q��?             B@������������������������       �������?             B@������������������������       �        `             c@w      �                   �?��j�`a�?�           d�@x                          �? �L�T�?{           @�@y      |                   �? >RR��?$           �{@z      {                   �?��e��?�            Pq@������������������������       �r�q��?             (@������������������������       � �Zz�q�?�            �p@}      ~                   �?�vPy`�?e            �d@������������������������       ��<ݚ�?             "@������������������������       ���e3���?`            �c@�      �                   �?�k2w��?W           `�@�      �                   �?t��}��?�            px@������������������������       ��n_Y�K�?             *@������������������������       �d�;lr�?�            �w@�      �                   �?�C��2(�?i            �d@������������������������       �      �?              @������������������������       ��f���?e            �c@�      �                    �?���%y�?c           ��@�      �                   �?��1G�v�?�             j@������������������������       �R���Q�?g             d@������������������������       �     ��?!             H@�      �                   �?�|�?�            v@������������������������       �f�n��,�?�            0r@������������������������       ��^�����?+             O@�      �                    �?P�x���?�           �@�      �                   �?�(\��e�?.            �@�      �                   �?0��:�*�?w           H�@�      �                   �?%}�p��?c             b@������������������������       �"pc�
�?             6@������������������������       �����v��?S            �^@������������������������       �h�v��+�?           ��@�      �                   �?��r
'��?�            pq@�      �                   �?և���X�?             E@������������������������       �                     @������������������������       �      �?             B@������������������������       � �\���?�            �m@�      �                   �?�dMƏ�?�           ,�@�      �                   �?��d~w�?           ��@�      �                   �?p�9�A��?�            @j@������������������������       ���p\�?            �D@������������������������       �X��ݥ��?l             e@������������������������       �p �_�G�?�           x�@�      �                   �?X��L���?           �y@�      �                   �?V{q֛w�?)             O@������������������������       ��q�q�?             @������������������������       �>4և���?$             L@������������������������       �81��=�?�            �u@�      �                   �?`*DB�?9           �@�      �                   �?$�,Y�&�?�           ̜@�      �                    �?v����?�           ��@�      �                   �?���eo�?�            @l@�      �                   �?H�U?B�?5            �T@������������������������       �                     "@�      �                   �?�1��u�?/            @R@������������������������       ��θ�?             :@������������������������       �                    �G@�      �                   �?tk~X���?^             b@������������������������       �h�����?J             \@������������������������       �      �?             @@�      �                   �?���aA�?           �{@�      �                   �?�6,r➷?�            �t@������������������������       �H%u��?             9@�      �                   �?�q���?�            s@������������������������       �����?'            @P@������������������������       �x�G�z�?�             n@�      �                   �?�h����?E             \@������������������������       �@3����?             K@������������������������       � _�@�Y�?'             M@�      �                   �?�g0�?�           \�@�      �                   �?t�BG_��?@           `�@�      �                   �?V�a�� �?             =@�      �                    �?�eP*L��?             &@������������������������       �X�<ݚ�?             "@������������������������       �                      @������������������������       �                     2@�      �                   �?�xO��?-           �~@�      �                    �? �g�oF�?�            pw@������������������������       ���Y��]�?e            �d@������������������������       ��S	���?z            `j@�      �                    �?�*;L�?N             ^@������������������������       ��θ�?)            @P@������������������������       ����Q��?%            �K@�      �                    �?:��V�?�           X�@�      �                   �?v�~��l�?�            @q@�      �                   �?�t����?             1@������������������������       �                     �?������������������������       �      �?             0@�      �                   �?+����?�            0p@������������������������       ��A�D6h�?g            �d@������������������������       �      �?B             W@�      �                   �?��xd�?�            pw@�      �                   �?�r����?            �F@������������������������       �      �?              @������������������������       �                    �B@�      �                   �?�'�`d�?�            �t@������������������������       ��!���?�            �m@������������������������       �JJ����?8            �W@�      �                    �? dB�?�           ݳ@�      �                   �?Ȟ�b׿?�           $�@�      �                   �?������?m           ��@�      �                   �?P����?K            �]@������������������������       �                     @������������������������       ��h����?F             \@������������������������       ��P)em�?"           �{@�      �                   �?����@��?           X�@�      �                   �?`�Q��?�             i@������������������������       ����N8�?/            �O@������������������������       ��z�>#h�?X             a@�      �                   �?�e<3��?�           8�@�      �                   �?����p�?�             q@������������������������       �                     �?������������������������       �0M����?�            �p@������������������������       ��#h���?�           ��@�      �                   �?P,9�u�?!           ��@�      �                   �?�#�˺�?�           ��@������������������������       �                    �E@�      �                   �?�U�:��?�           H�@�      �                   �?J�yE�?�            �o@������������������������       � pƵHP�?a            �c@������������������������       �X&$�E�?@            �X@������������������������       �8��㋱?           �x@�      �                   �?Xs�' ��?g           @�@������������������������       � $����?}           ȏ@�      �                   �?�#-���?�           ��@������������������������       �R�vz ��?�            �h@������������������������       ��-T�J�?j           ��@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B0      �h�@    ���@     ��@     X�@    ���@      �@     T�@     X�@     �@     �{@     �@     �{@     �z@     �r@     �z@     �r@      l@     `h@     `i@      Z@      �?             �S@      b@     @S@      b@      �?                       @     ��@     �v@     P�@     �b@     �a@      @     �Z@      @     �Z@       @      V@       @      3@                      �?     �@@       @      =@      �?      @      �?      �@      b@     P�@     �P@     �@      H@     ��@      B@     ��@      ?@     8�@      >@      8@      �?     pu@      @     �s@      @      ?@             �F@      (@     �D@      (@      @              @      3@       @      (@      @      @      @      @      �?       @     �u@     �S@     @t@      G@     �i@     �E@     �i@      B@     `h@     �A@      &@      �?      �?      @     @]@      @     @]@      �?     �X@      �?      3@                       @      :@      @@      :@      9@      4@      9@      @                      @     �q@     �j@     �q@     @e@     Pp@      `@      c@     @V@     �Z@     �D@     �Y@      B@      @      @      G@      H@      E@      H@      @              [@      D@     �W@      B@      R@      1@      6@      3@      ,@      @      @       @      "@       @      7@     �D@      ,@      7@      "@      2@      @      2@      @                     �F@    �\�@     T�@    ���@     @y@     ��@      v@     l�@     `h@     x�@      4@     �@      3@     ��@      "@      Z@             �@      "@     H�@      $@      ,@             ؃@      $@     �@      �?      K@             8�@      �?     ��@             �~@      �?     `�@     �e@     �@     �Y@     t�@      O@      @             h�@      O@     ��@      D@      �?             ��@      D@     ��@     @R@     �@      ?@      @             ؄@      ?@     (�@      E@      @              �@      E@     ��@     �c@     P�@      &@     ��@      $@     �u@      @      o@      @     �w@      �?     �k@      �?     `c@             (�@     @b@     ��@     @R@     �z@     �C@     �|@      A@     ��@     @R@     s@     �G@     �l@      :@     ܐ@      J@     ��@      A@     �r@      �?      @             �r@      �?     �g@      �?     �Z@             0{@     �@@     �m@      1@     �h@      0@     �u@      2@      Z@      �?     �N@             �E@      �?      n@      1@     `a@      ,@     �Y@      @     �@     �@     ȇ@     `s@     �x@     �b@     �n@     �X@      c@      I@     �v@     @d@     �p@      _@      c@     �T@     �\@      E@      X@      C@      K@      1@      E@      5@     �|@     �t@     `v@      q@     @i@      d@     �Z@     @T@      X@     �S@     �c@     �\@      Y@     �Q@      L@     �E@     �X@     �L@     �H@      <@      I@      =@     h�@     �@     �u@     8�@      k@     $�@     �]@     Px@              �?     �]@     @x@     �W@     Pu@      &@     �e@      &@     �`@             �D@     �T@      e@      I@     �Y@     �@@     �P@      9@     �G@      "@      7@      0@      8@     @X@      �@     @R@     x�@     �F@     �v@      <@      l@      8@     @]@     �`@     (�@     @\@      �@      S@     P|@      @      `@              @      @     �^@      R@     @t@     �C@      Q@     �@@      p@               @     �@@     �o@     �B@     `k@              �?     �B@     @k@      =@     �Q@      �?      D@      <@      ?@       @     `b@      5@     �l@              �?      5@     �l@      *@      U@       @      I@      &@      A@       @      b@     �m@     ��@     `f@     ��@     �\@     \�@     @Q@     �@             �b@     @Q@     `�@     �D@     �T@      <@     �{@     �F@     ��@      @      `@      E@     @@      2@     �Q@      8@     �z@     @P@     h�@     �E@     Pr@      =@     @Y@              M@      =@     �E@      ,@      h@      6@     �r@              E@      6@     �o@      @      <@      1@     @l@      N@     0�@      <@      l@      *@     �^@      �?      U@      (@     �C@      .@     �Y@      @      O@      (@      D@      @@     (�@      0@     �l@      0@     r@     �@     ��@     A�@    �G�@     x�@     ��@     t�@     �@     ؜@     `v@     Ȓ@     s@     �\@      m@      @     @V@      @      *@      �?      S@     �Z@     �a@      H@     �M@      B@     �M@      (@             �M@      U@     �K@      U@      @              �@     @R@     �v@      @     @g@      @      @             �f@      @      f@      @      �?              f@      @     ��@     �P@     �v@      =@     �v@     �B@      �@     �J@     �k@     �@@     ``@      &@      @      �?      �?      �?       @              `@      $@      D@      $@      V@              W@      6@      ,@      5@              �?      ,@      4@     �S@      �?      �?             @S@      �?     Pz@      4@     �j@      ,@      @             @j@      ,@     �i@      @      @             �i@      @     @p@     �f@      g@     @_@     �R@     �Q@      �?      8@     @R@      G@     �[@     �K@       @      *@      [@      E@      S@      M@      G@     �@@              @      G@      ;@      >@      9@              @      >@      3@      p@     �@      "@     h�@       @     @m@      �?     �g@              4@      �?      e@      �?     �F@              @      �?      E@      @     0z@      @     �u@             �R@      @     q@       @      R@      o@     ��@     `b@     Pp@     @P@      ]@     �E@     �R@      6@     �D@     �T@      b@     �Q@     �Z@      &@     �C@     �Y@     ��@      P@      �@     �G@     u@              �?     �G@      u@      1@     0{@              @      1@     �z@      C@     @r@      0@     �a@      6@     �b@     �@     ��@     T�@     :�@      x@     .�@      g@     8�@      g@     �j@     �_@     �g@      7@     �f@      Z@      @     �L@      :@       @      8@     �K@       @             ��@     @i@     ��@      d@     �@     �c@     �}@      7@     P}@      a@      @       @     ��@     �D@     �f@     �D@      ?@      @      >@     �A@      �?              c@     L�@     0�@      �@     �`@     �x@      G@     �n@     �@@      $@       @     @m@      ?@     @c@      *@      @       @     `b@      &@     `}@     �U@      t@     �Q@       @      @     �s@     �P@     �b@      .@      @      �?     �a@      ,@     �e@      x@     �L@     �b@      B@      _@      5@      ;@     �]@     `m@     @V@     @i@      =@     �@@      w@     6�@     �c@     ��@     �_@     X�@      Q@     @S@      @      2@      P@     �M@      M@     ��@      >@      o@      2@      8@              @      2@      2@      (@      l@     �j@     ܘ@     `d@     4�@      Z@     �Z@      @      C@     @Y@      Q@     �M@     ��@     �H@     �v@      ;@     �A@      @       @      7@     �@@      6@     pt@     Ė@     _�@     ܑ@     ��@     �j@     `|@      V@     @a@     �J@      =@              "@     �J@      4@      @      4@     �G@             �A@     @[@      @      [@      ?@      �?     �_@     �s@      0@     �s@      @      6@      *@     @r@      @     �N@      "@     �l@     �[@       @     �J@      �?     �L@      �?     �@     �n@     �{@     �T@      @      7@      @      @      @      @       @                      2@     @{@     �M@     v@      6@      d@      @      h@      2@     �T@     �B@      I@      .@     �@@      6@     p~@     �d@     �k@     �K@       @      .@      �?              �?      .@     `k@      D@     �b@      1@     @Q@      7@     �p@     @[@      @     �C@      @       @             �B@     @p@     �Q@     @j@      :@      I@      F@     �s@     ��@      ^@     D�@      @     p�@       @      ]@              @       @     �[@      @     �{@     �\@     ��@      P@      a@      .@      H@     �H@      V@     �I@     ؎@      4@     �o@              �?      4@     `o@      ?@     ��@     @h@     $�@     �K@     �@             �E@     �K@     ��@     �D@     �j@      @      c@      C@     �N@      ,@     �w@     `a@     *�@      @     ��@     �`@     ��@     �P@     �`@      Q@     p�@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h7Kh8Kh9h"h#K �r�  h%�r�  Rr�  (KK�r�  hQ�C              �?r�  tr�  bhEhUh@C       r�  �r�  Rr�  hYKhZh[Kh"h#K �r�  h%�r�  Rr�  (KK�r�  h@�C       r�  tr�  bK�r�  Rr�  }r�  (hKheM�hfh"h#K �r�  h%�r�  Rr�  (KM��r�  hm�B�e                             �?��6��?�e           �@       �                    �?*Zfa��?�4          ��@       d                    �?�&ӿ��?x(          ��@       I                    �?=
M1%�?�          ���@                            �?(8�O�?p           ��@������������������������       �ܤm6��?           �y@       .                    �?����i/�?j           ��@                           �?��;�;j�?3           ��@	                           �?ʽ�C�?�           ��@
                            �?�p ��?I           ��@������������������������       ��q@{)�?�            �q@������������������������       �T�7�4�?�             o@                           �?�d	���?f            �c@                            �?�f���?e            �c@                           �?��x$�?I            �\@                           �? T���v�?H            @\@������������������������       �г�wY;�?@            �Y@������������������������       �                     &@������������������������       �                      @                           �?0,Tg��?             E@                           �?�E��ӭ�?             B@������������������������       ��t����?             A@������������������������       �                      @������������������������       �r�q��?             @������������������������       �                     �?       %                     �?�ep���?�           x�@                           �?�`>:��?�           ,�@������������������������       �                     @       "                    �?�0���?~           �@       !                    �?h�=V��?R           (�@                            �?p�u$v��?1           H�@������������������������       ��č����?v           ��@������������������������       �H��M��?�            �r@������������������������       ��������?!             N@#       $                    �?Pa�	�?,            �P@������������������������       ��C��2(�?             6@������������������������       �                     F@&       +                    �?V6q�_�?           0y@'       *                    �?H�o����?�            @w@(       )                    �?K�� ��?�            `u@������������������������       ��n����?�            �m@������������������������       ��&=�w��?D            �Z@������������������������       ���S���?             >@,       -                    �?��a�n`�?             ?@������������������������       �@�0�!��?	             1@������������������������       �                     ,@/       <                     �?P�(�&b�?7          ���@0       1                    �?`��o�?-           [�@������������������������       �        ^            ``@2       7                    �?0!�����?�           ص@3       6                    �?�/��l�z?�           z�@4       5                    �? N�Tov?Y           �@������������������������       ��,X����?k           ��@������������������������       �        �           H�@������������������������       � �ׁsF�?w             i@8       9                    �?\��A��?�           6�@������������������������       �hY����?�           ��@:       ;                    �?�y�9&/�?           ؙ@������������������������       ��V����?S           ؔ@������������������������       �     �?�             t@=       >                    �?�6�Z�5�?
           ��@������������������������       �                    �H@?       D                    �?`�5
��?�           6�@@       A                    �?�H���?           |�@������������������������       � �,�:�?�           ��@B       C                    �?�^��3|?q           �@������������������������       ����C-��?>           �~@������������������������       �        3            �U@E       F                    �?�#�S�`�?�           �@������������������������       ����y�?�           ��@G       H                    �? \sF��?7           @�@������������������������       ����7�?�            �@������������������������       �`2U0*��?|             i@J       S                    �?4�W��?3           ��@K       N                     �?�so=���?=           �@L       M                    �?x�dPS[�?�            pq@������������������������       ��t`�4 �?R            �^@������������������������       ��*���^�?`            �c@O       P                    �?�l�Z-��?�            `l@������������������������       �                     @Q       R                    �?6���?�            �k@������������������������       ��KM�]�?=            �W@������������������������       �tϺFˁ�?J            @_@T       ]                    �?�-����?�            Px@U       X                     �?xdQ�m��?d            @d@V       W                    �?��y� �?6            @W@������������������������       �                    �F@������������������������       �r�q��?             H@Y       \                    �?��.N"Ҭ?.            @Q@Z       [                    �?�?�|�?            �B@������������������������       �                      @������������������������       ���?^�k�?            �A@������������������������       �      �?             @@^       a                    �?^��8g�?�            `l@_       `                     �?��S���?b            �b@������������������������       ��eP*L��?:             V@������������������������       ��g�y��?(             O@b       c                     �?���|���?0            @S@������������������������       �������?            �D@������������������������       �X�<ݚ�?             B@e       �                    �?��=���?�
            �@f       �                    �?�������?.           Ʃ@g       x                    �?���~e��?�           С@h       m                    �?�̗����?&           P}@i       j                     �?@�r-��?F            �]@������������������������       �և���X�?            �A@k       l                    �?P��BNֱ?3            �T@������������������������       �Ћ����?2            �T@������������������������       �                     �?n       s                     �?z�����?�            �u@o       r                    �?>4և���?k             e@p       q                    �?Rg��J��?^            `b@������������������������       �ؓ��M{�?G            �[@������������������������       ���G���?            �B@������������������������       �                     5@t       w                    �?�n/S��?u            �f@u       v                    �?<=�,S��?o            �e@������������������������       �ꟲ�4��?X            @a@������������������������       ���+��?            �B@������������������������       �                      @y       �                     �?n��r�?v           L�@z                           �?p��l?�?N           Ќ@{       |                    �?�tVV�?f           ��@������������������������       �                     @}       ~                    �?h]���~�?d           ��@������������������������       ��˫���?y             g@������������������������       �P��a4�?�            �w@�       �                    �?�-��?�            `v@������������������������       �                     @�       �                    �?�Yre��?�             v@������������������������       �        C             Z@������������������������       �ףp=
�?�            @o@�       �                    �?��O*��?(           ȋ@������������������������       �                     @�       �                    �?��@���?%           ��@�       �                    �?8:U��ܻ?~           ��@������������������������       �XB���?u            `i@������������������������       �������?	           0y@�       �                    �?��?^�k�?�            �q@������������������������       ��?�|�?/            �R@������������������������       � f^8���?x            �i@�       �                    �?&�Z���?�           ؏@�       �                    �?�|\Ur�?            ؈@�       �                    �?     ��?M            �@������������������������       �        6            �T@�       �                     �?0!kp���?           �z@������������������������       �@ o����?k            �d@������������������������       ��X�G�U�?�            �p@�       �                     �?\m�����?�            �q@������������������������       �l��
I��?A             [@������������������������       �]�	�?r            �e@�       �                    �?     ��?�             l@������������������������       �                     �?�       �                    �?t�R2��?�            �k@�       �                     �?��:�-�?D            @Y@������������������������       ���<b�ƥ?             G@������������������������       � �Jj�G�?&            �K@�       �                     �?����5�?M            �^@������������������������       �V��z4�?%             O@������������������������       ���Q��?(             N@�       �                    �?��d��?�           ��@�       �                    �?^(��I�?s           �@�       �                     �?��"Ҥ(�?U            �b@�       �                    �?��|�5��?            �G@������������������������       �                      @�       �                    �?��Hg���?            �F@������������������������       ��KM�]�?             C@������������������������       �                     @�       �                    �?$�q-�?:             Z@������������������������       �                    �@@�       �                    �?�Z��L��?)            �Q@������������������������       ���ɉ�?'            @P@������������������������       �                     @�       �                     �?�D�n���?           `|@�       �                    �?0��X�t�?|            �h@������������������������       �                    �H@������������������������       ���<�Ұ?^            `b@�       �                    �?֨!t��?�             p@������������������������       ��&=�w��?            �J@������������������������       ���p\�?�            �i@�       �                    �?p=
ף0�?4            ~@������������������������       �                    �C@�       �                     �?؇���X�?           �{@�       �                    �?�R����?n            �e@������������������������       ���:�-�?A            @Y@������������������������       �ޚ)�?-             R@�       �                    �?��v����?�            �p@������������������������       ��B:�g�?t            �e@������������������������       ����!���?<            �W@�       �                    �?��d?S��?s           ��@�       �                    �?\u�S>�?L           �@�       �                     �?�7��d��?A             Y@�       �                    �?�����H�?            �F@�       �                    �?�S����?             3@�       �                    �?@4և���?
             ,@������������������������       ��C��2(�?             &@������������������������       �                     @������������������������       ����Q��?             @�       �                    �?$�q-�?             :@������������������������       �r�q��?             (@������������������������       �        	             ,@�       �                    �?h㱪��?#            �K@�       �                    �?�IєX�?             1@������������������������       ��8��8��?             (@������������������������       �                     @�       �                    �?P�Lt�<�?             C@������������������������       �P���Q�?             4@������������������������       �                     2@�       �                    �?�р�q�?           X�@�       �                     �?����b�?           8�@�       �                    �?DheST��?            {@������������������������       �����X�?�            �t@������������������������       �$+ޠ�5�?H            @Z@�       �                    �?��
���?�            Pw@������������������������       �:��Z��?�            @k@������������������������       ��@1B�?_            `c@�       �                     �?j����?           x�@�       �                    �?b�'����?!           �|@�       �                    �?�/C��?�            �t@������������������������       ��
�G�?�            �p@������������������������       ���M��?.            �Q@�       �                    �?d58��1�?N            �^@������������������������       �д>��C�?&             M@������������������������       �     ��?(             P@�       �                    �?p�����?�            `v@�       �                    �?�1��u�?�            `k@������������������������       ��J�j�?e            �c@������������������������       �ƆQ����?(            �N@�       �                    �?t�0i��?W            `a@������������������������       ���&����?&            @P@������������������������       ��Gi����?1            �R@�       �                    �?4,Y$�?'           ��@������������������������       �                     4@�       �                    �?�ȡp�(�?           b�@�       �                     �?���Ĩ��?�           Ģ@�       �                    �?ДX��?           0�@�       �                    �?�<����?�           0�@������������������������       �/�%��?            0z@������������������������       ����f\1�?�            0z@�       �                    �?`BP���?           `|@������������������������       �l�?����?�            �q@������������������������       ��}�+r��?g            `e@�       �                    �?�j�LD�?�           X�@�       �                    �?d�S����?�           h�@������������������������       ��l�ո�?�            `r@������������������������       ����_�?           p|@�       �                    �?������?�            �v@������������������������       ��8��8��?q             h@������������������������       �$�Q�\�?h             e@�       �                     �?���:b�?i           x�@�       �                    �?�S���?           �y@������������������������       �4��?�?a            �c@������������������������       �@���|N�?�             p@�       �                    �?��6��?b           ��@������������������������       � d��u�?R            @_@������������������������       ��~�y�C�?           @{@      f                   �?_	�?�0          �.�@      E                   �? U�<��?�           ۻ@      2                   �?�@�;���?m
           C�@                         �?������?�           ��@                         �?"�s%��?           ̟@                         �?�ᨰ�l�?1           �@      
                    �?�wV����?#           X�@      	                   �?��4�&��?H           ��@������������������������       �^Z�sl�?b            �b@������������������������       � n<�(�?�            �w@                         �?�߄��?�            �u@                         �?�p ��?3            �T@������������������������       �      �?              @������������������������       �z�G���?1             T@������������������������       �����e��?�            �p@                         �?�y+v�?           p�@                          �?؇���X�?             5@������������������������       �"pc�
�?             &@������������������������       �ףp=
�?             $@                          �?�M)��?           ȇ@������������������������       �(;�ŀ	�?2           @|@������������������������       �\�t��Y�?�            Ps@                         �?�p�Ү��?�            �w@������������������������       �                     6@                          �?r�����?�            @v@������������������������       ���V�j��?z            �h@������������������������       ������?c            �c@      '                   �?�#k~��?�           P�@      "                    �?p�|����?O            @\@      !                   �?�d�����?4             S@                          �?��X���?/            @Q@������������������������       ���f/w�?)            �N@������������������������       �                      @������������������������       �                     @#      &                   �?؀�:M�?            �B@$      %                   �?V�a�� �?             =@������������������������       �      �?             8@������������������������       �                     @������������������������       �                      @(      /                   �?�
l?�?]           ��@)      ,                   �?��&�J޸?�           ��@*      +                    �? ���l�?�            @x@������������������������       � "���?�            pp@������������������������       �@�n�1�?Y            @_@-      .                    �?�m�&��?�           H�@������������������������       ��l�+���?           P}@������������������������       �p��%���?�            @q@0      1                    �?4\O�ޕ�?�            �n@������������������������       ��G�z��?a             d@������������������������       �h�|�`�?7            �U@3      :                   �? 9��w��?�           ��@4      9                   �?V�a�� �?8            �U@5      8                   �?�+e�X�?2            �R@6      7                    �?��oh���?0            @R@������������������������       ��d�����?             C@������������������������       �b�h�d.�?            �A@������������������������       �                      @������������������������       �                     (@;      @                    �?��K#u��?l           (�@<      ?                   �?�N5X��?�            r@=      >                   �?h��)�~�?�            @l@������������������������       �����e��?-            �P@������������������������       �p=
ף0�?e             d@������������������������       �b����?-            �O@A      D                   �?�?�<��?�            @p@B      C                   �?x�û��?w             g@������������������������       �0�,���?'            �P@������������������������       �@\�*��?P            @]@������������������������       ����=A�?6             S@F      O                   �?�s��=�?O           0�@G      J                    �?0�����?f           ��@H      I                   �?@ux�ᭉ?�            �s@������������������������       ��NM�g�?a            �e@������������������������       �        X             b@K      L                   �?��.N"Ҭ?�            @q@������������������������       �`'�J�?`             c@M      N                   �?�-.�1a�?M            �^@������������������������       �                     I@������������������������       ���pBI�?.            @R@P      [                   �?��D×
�?�           ��@Q      V                    �?�f��9��?#           0}@R      U                   �?����,�?�            @q@S      T                   �?��_����?�            �k@������������������������       ����@M^�?O             _@������������������������       ����Q �?7            �X@������������������������       ��E��ӭ�?              K@W      X                   �?����%��?}            �g@������������������������       �� ���?A            @Z@Y      Z                   �?"Z�l�?<            �U@������������������������       ���hJ,�?             A@������������������������       �8�Z$���?$             J@\      _                   �?D���D|�?�           Н@]      ^                    �?�ہ��?K           ��@������������������������       ������?3           �}@������������������������       ��\|X��?           P|@`      c                   �?�����?{           ��@a      b                    �?\ ���?.           �}@������������������������       �8���@�?�            `m@������������������������       �H�4�l��?�            �m@d      e                    �?������?M           �@������������������������       �8��?�A�?�             k@������������������������       �h�a��?�            0r@g      �                   �?��3u�'�?�          �o�@h                         �?8��x���?�           �@i      t                    �?����'2�?7           �@j      o                   �?��P���?�           x�@k      n                   �?�Q���J�?Z           `�@l      m                   �?$���s�?�            Pu@������������������������       �T��mh��?�             l@������������������������       ����"�?H             ]@������������������������       � :�|Nk?w           ��@p      s                   �?\{��)x�?m            @f@q      r                   �?ƈ�VM�?4            @V@������������������������       �z�G�z�?            �F@������������������������       �`���i��?             F@������������������������       �        9            @V@u      |                   �?`�AזI�?p           h�@v      y                   �?�S{��?�           �@w      x                   �?FH5�j�?h           ��@������������������������       �H� >ſ�?           |@������������������������       �h�����?I             \@z      {                   �?#z�i��?/            �T@������������������������       ��4F����?            �D@������������������������       �                    �D@}      ~                   �? ��t?�           \�@������������������������       � Mk�9�n?�           ��@������������������������       � �w5�?K            �]@�      �                    �?����ź?�           �@�      �                   �?��"�?k           ��@�      �                   �?�Y�R_�?\            �a@������������������������       �0��_��?E            �Z@������������������������       ��X�<ݺ?             B@������������������������       � �0�G�r?            {@�      �                   �?�J�
;�?O           ��@�      �                   �?�Y�����?�            �s@������������������������       �\����?�            pp@������������������������       ��1�`jg�?'            �K@������������������������       �        �           ��@�      �                    �?vE�*4��?           �@�      �                   �?T�����?�           ��@�      �                   �?~$�����?n           ؎@�      �                   �?:tl3.��?           �{@�      �                   �?�����?�            �q@������������������������       ��q�q�?             @������������������������       �H�_��?�            0q@������������������������       �"�W1��?m            �d@�      �                   �?��R(�<�?W           ��@�      �                   �?������?�            @k@�      �                   �?=0�_�?]             c@������������������������       �؇���X�?             @������������������������       ��c!�^�?W            @b@������������������������       ��	j*D�?&            @P@�      �                   �?\AUj��?�            @t@�      �                   �?p^�AL�?{            �g@������������������������       �                      @������������������������       ������H�?y            �g@������������������������       ������B�?Y            �`@�      �                   �?L��JT�?           �@�      �                   �?�;���?           ܒ@�      �                   �?@��T�?[           P�@�      �                   �?��S���?\            �`@������������������������       �H%u��?             9@������������������������       ��eP*L��?N            �[@������������������������       �@k��s�?�           �@�      �                   �?�:c�t�?�            �p@�      �                   �?��c:�?             G@������������������������       �                     @������������������������       ��lg����?            �E@������������������������       �������?�            �k@�      �                   �?�%���?           P�@�      �                   �?+Y���?G            @\@������������������������       ��8��8��?             8@������������������������       �����?9            @V@������������������������       � k_��?�           Ȇ@�      �                   �?�V���?|           �@�      �                   �?෹�A��?9           ��@�      �                   �?ȼ�F��?�            �@�      �                   �?<���D�?            �@@�      �                   �?���y4F�?             3@������������������������       �      �?	             (@������������������������       �؇���X�?             @������������������������       �                     ,@�      �                   �?�[d"(�?�           �@������������������������       ��S3��?�             t@�      �                   �?`�ǆ�3�?           z@������������������������       ��h�*$��?e             c@������������������������       �̘#ZJ�?�            �p@�      �                   �?��4ȅ�?M           ��@������������������������       �θ	j*�?�            @p@�      �                   �?��1|���?�            �q@������������������������       ��b��[��?'            �K@������������������������       �P����?�            �l@�      �                   �?LLڥ=��?C           ک@�      �                   �?      �?�            �w@�      �                   �? ,U,?��?3            �T@�      �                   �? i���t�?            �H@������������������������       �`Ӹ����?            �F@������������������������       �      �?             @������������������������       �                     A@�      �                   �?>�O��?�            �r@�      �                   �?�1׹k��?�            �h@������������������������       �F��U@�?g            @c@������������������������       �X��ʑ��?            �E@������������������������       ��\�u��?<            �Y@�      �                   �?HI��ڻ?R           ަ@������������������������       ����̺��?�           �@�      �                   �?hSA�k�?S           ��@������������������������       ��FVQ&�?�            �t@������������������������       � kV�X�?n           |�@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KM�KK�r�  hQ�B      �l�@    ���@    �m�@     S�@     ��@     ��@     ��@     ��@     �@     ��@     �i@     @i@     ��@     `�@     ��@     �z@     0y@      r@     @p@     q@     �d@     �]@     �W@     @c@     �a@      .@     �a@      ,@      \@      @     �[@      @     �X@      @      &@               @              ?@      &@      :@      $@      8@      $@       @              @      �?              �?     X�@      a@     H�@     �P@      @             (�@     �P@     (�@      P@     ��@      I@     ��@      D@     r@      $@      G@      ,@      P@       @      4@       @      F@             �t@     �Q@     s@     �P@     r@     �J@     `g@     �H@     �Y@      @      0@      ,@      <@      @      ,@      @      ,@            �a�@     �l@     ϵ@     �a@     ``@             L�@     �a@     h�@      "@     ܣ@      @     p�@      @     H�@             �h@       @     0�@     ``@     ��@     �O@     Ș@      Q@     �@     �J@     s@      .@     �@      V@     �H@             ��@      V@     \�@       @     ��@      @     �@       @     �~@       @     �U@             ��@      T@     `�@      D@      �@      D@      �@      @@      h@       @     @m@     ��@     �_@     �w@     �P@     �j@      &@     �[@      L@     @Y@     �M@      e@              @     �M@      d@      $@     @U@     �H@      S@      [@     �q@      $@      c@       @     @U@             �F@       @      D@       @     �P@      �?      B@               @      �?      A@      �?      ?@     �X@      `@     �Q@      T@      D@      H@      >@      @@      <@     �H@      (@      =@      0@      4@      �@     @�@     �@     T�@     ȝ@     `w@     �g@     pq@      2@      Y@      .@      4@      @      T@      @     �S@              �?     �e@     `f@     �X@     @Q@     �S@     @Q@      H@      O@      >@      @      5@             @R@     �[@     @P@     �[@     �G@     �V@      2@      3@       @             К@     �W@     0�@      J@     Ȁ@      ;@      @             ��@      ;@     `f@      @      v@      6@     �t@      9@      @             �t@      9@      Z@              l@      9@     p�@     �E@      @             X�@     �E@     ؁@     �A@     �h@      @     pw@      <@      q@       @      R@       @      i@      @     �c@     ��@     �\@     H�@      "@     p@             �T@      "@     Pz@       @     `d@      @      p@     @Z@     @f@      @@      S@     @R@     �Y@      E@     �f@              �?      E@     �f@       @     �X@      �?     �F@      �?      K@      D@     �T@      3@     �E@      5@     �C@     �@     ؁@     0|@     @c@      3@     �`@      &@      B@               @      &@      A@      @      A@      @               @      X@             �@@       @     �O@       @     �O@      @              {@      6@     �g@      @     �H@             �a@      @      n@      1@     �I@       @     �g@      .@     �O@     z@             �C@     �O@     �w@      ;@     @b@       @     �X@      9@     �G@      B@      m@      �?     �e@     �A@     �M@     ��@     ��@     �@     ��@      @     @W@      @      D@      @      0@      �?      *@      �?      $@              @       @      @       @      8@       @      $@              ,@       @     �J@      �?      0@      �?      &@              @      �?     �B@      �?      3@              2@     ��@     �}@     �@     �l@     �r@     ``@     `m@     �W@      Q@     �B@      q@     �X@     @e@      H@      Z@     �I@     ��@     `n@     t@      a@     �l@     �Z@      f@     �U@     �I@      4@     @W@      =@      H@      $@     �F@      3@     `o@     �Z@     �c@      N@      \@      G@     �G@      ,@      W@     �G@      H@      1@      F@      >@     0r@     D�@              4@     0r@     �@      l@     �@     �`@     �@      W@     P�@     �B@     �w@     �K@     �v@     �D@     �y@      @@     `o@      "@     @d@     �V@     ؏@     �L@     ��@     �D@     �o@      0@     p{@      A@     pt@      0@      f@      2@     �b@     �P@     `�@     �A@     �w@      .@     �a@      4@     �m@      @@     ��@      ,@     �[@      2@      z@     ׸@    ���@     B�@     t�@     $�@     ��@     N�@      �@     p�@     pu@      �@      f@     `�@     �W@      ~@     �H@     @[@     �D@     0w@       @     �r@      G@      D@      E@      �?      �?     �C@     �D@     @p@      @     ��@     �T@      2@      @      "@       @      "@      �?     P�@     �S@     �y@     �E@     q@      B@     �j@     �d@              6@     �j@      b@     @[@     @V@     �Y@     �K@     ,�@      i@     �S@      A@      L@      4@      L@      *@      H@      *@       @                      @      7@      ,@      7@      @      2@      @      @                       @     �@     �d@     ̐@      M@     x@      @     `p@      �?     �^@       @     ��@     �K@     �z@     �C@     @p@      0@      a@     @[@      V@      R@     �H@     �B@     �~@      b@      2@     @Q@      2@     �L@      0@     �L@      $@      <@      @      =@       @                      (@     �}@      S@     �n@      F@     �i@      6@     @P@      �?     `a@      5@     �D@      6@     �l@      @@      f@      @     @P@       @      \@      @     �I@      9@     �p@     �@      $@     8�@       @     �s@       @     `e@              b@       @     �p@      @     `b@       @     @^@              I@       @     �Q@     Pp@     ��@      `@      u@     @X@     `f@     �T@     �a@      H@      S@      A@      P@      .@     �C@      @@     �c@      3@     �U@      *@     @R@      @      =@       @      F@     �`@     ��@      K@     @�@      <@     �{@      :@     �z@     �S@     @�@      D@      {@      3@      k@      5@     @k@      C@     `}@      7@     @h@      .@     @q@     l�@    �T�@     �}@     �@      w@     �@     @g@      �@     �`@     0�@     �`@      j@      6@     `i@     �[@      @      �?     ��@      J@     �_@      J@     �B@      "@      B@     �E@      �?             @V@      g@     ��@     �f@     �|@     �_@      {@      3@     �z@      [@      @      K@      <@      *@      <@     �D@              @     P�@       @     |�@      �?     @]@     �Z@     D�@     �F@     ��@      F@     �X@      $@      X@      A@       @      �?     �z@     �N@      �@     �N@     p@      "@     �o@      J@      @             ��@     ��@     ��@     ��@     ��@     ��@     �s@     �q@     `d@      o@     �@@      @       @     �n@      ?@      A@     @`@      x@     �c@     �d@     �J@      b@       @      @      �?     `a@      @      4@     �F@     �k@     �Y@     @e@      5@       @              e@      5@     �I@     �T@      o@      �@      d@     X�@     �\@     ��@     �O@      R@      @      6@      N@      I@     �I@     ��@     �G@     �k@      ;@      3@              @      ;@      0@      4@     `i@      V@     ��@      N@     �J@       @      6@      M@      ?@      <@     �@     �@     ��@     �@     `|@     8�@     @W@      =@      @      .@      @      "@      @      @      �?      ,@             P�@     @V@     �p@     �I@     �w@      C@      a@      .@     @n@      7@     �f@     �v@     @U@     �e@     @X@     @g@      3@      B@     �S@     �b@     �v@     
�@     �g@     �g@      @     �S@      @      F@       @     �E@      @      �?              A@     @g@     @\@      ]@     @T@     �W@     �M@      5@      6@     �Q@      @@      e@     ��@      O@      �@     �Z@     ��@      4@     `s@     �U@      �@r�  tr�  bubhhubehhub.